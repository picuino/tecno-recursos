CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
21 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
19
9 Resistor~
219 414 100 0 1 5
0 0
0
0 0 608 0
2 1k
-7 -14 7 -6
2 R5
-6 -12 8 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5993 0 0
2
44525.6 0
0
7 Ground~
168 390 210 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8654 0 0
2
44525.6 0
0
2 +V
167 419 190 0 1 3
0 5
0
0 0 53344 180
4 -15V
-13 12 15 20
2 V3
-5 0 9 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7223 0 0
2
44525.6 2
0
2 +V
167 419 132 0 1 3
0 6
0
0 0 53344 0
3 15V
-11 -27 10 -19
2 V4
-7 -15 7 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3641 0 0
2
44525.6 1
0
8 Op-Amp5~
219 419 159 0 5 11
0 2 4 6 5 3
0
0 0 64 0
5 UA741
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 1 0 0
1 U
3104 0 0
2
44525.6 0
0
9 Resistor~
219 339 185 0 1 5
0 0
0
0 0 608 0
2 1k
-7 -14 7 -6
2 R4
-6 -12 8 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3296 0 0
2
44525.6 0
0
9 Resistor~
219 338 153 0 1 5
0 0
0
0 0 608 0
2 1k
-7 -14 7 -6
2 R3
-6 -12 8 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 62
82 0 0 0 1 0 0 0
1 R
8534 0 0
2
44525.6 0
0
2 +V
167 269 186 0 1 3
0 5
0
0 0 53344 180
4 -15V
-13 12 15 20
2 V2
-5 0 9 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
949 0 0
2
44525.6 11
0
2 +V
167 269 126 0 1 3
0 6
0
0 0 53344 0
3 15V
-11 -27 10 -19
2 V1
-7 -15 7 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3371 0 0
2
44525.6 10
0
8 Op-Amp5~
219 269 153 0 5 11
0 2 4 6 5 3
0
0 0 64 0
5 UA741
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 1 0 0
1 U
7311 0 0
2
44525.6 9
0
7 Ground~
168 157 208 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3409 0 0
2
44525.6 8
0
10 Capacitor~
219 193 147 0 2 5
0 4 7
0
0 0 576 180
6 0.01uF
10 0 52 8
2 C1
-7 -18 7 -10
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3526 0 0
2
44525.6 7
0
11 Signal Gen~
195 47 152 0 64 64
0 8 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 18
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 64 0
5 -1/1V
-18 -30 17 -22
2 Vi
-6 -33 8 -25
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 1 0 0
1 V
4129 0 0
2
44525.6 6
0
7 Ground~
168 228 208 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6278 0 0
2
44525.6 5
0
7 Ground~
168 85 208 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3482 0 0
2
44525.6 4
0
10 Capacitor~
219 196 62 0 2 5
0 7 3
0
0 0 576 0
6 0.02uF
-22 -18 20 -10
2 C2
-6 -20 8 -12
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8323 0 0
2
44525.6 3
0
9 Resistor~
219 157 179 0 3 5
0 2 7 -1
0
0 0 608 90
2 1k
8 0 22 8
2 Rr
4 -7 18 1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3984 0 0
2
44525.6 2
0
9 Resistor~
219 267 91 0 2 5
0 4 3
0
0 0 608 0
6 11.25k
-21 -14 21 -6
2 R2
-5 -13 9 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7622 0 0
2
44525.6 1
0
9 Resistor~
219 128 147 0 2 5
0 8 7
0
0 0 608 0
6 11.25k
-21 -14 21 -6
2 R1
-4 -14 10 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
816 0 0
2
44525.6 0
0
22
5 2 0 0 0 0 0 5 1 0 0 4
437 159
461 159
461 100
432 100
0 1 0 0 0 0 0 0 1 4 0 3
373 153
373 100
396 100
1 1 0 0 0 0 0 2 5 0 0 3
390 204
390 165
401 165
2 0 0 0 0 0 0 6 0 0 5 3
357 185
373 185
373 153
2 2 0 0 0 0 0 7 5 0 0 2
356 153
401 153
1 4 5 0 0 0 0 3 5 0 0 2
419 175
419 172
1 3 6 0 0 0 0 4 5 0 0 2
419 141
419 146
1 0 0 0 0 0 0 6 0 0 21 5
321 185
303 185
303 232
102 232
102 147
1 0 0 0 0 0 0 7 0 0 19 2
320 153
303 153
1 1 2 0 0 0 0 10 14 0 0 3
251 159
228 159
228 202
2 0 3 0 0 0 0 18 0 0 19 2
285 91
303 91
1 0 4 0 0 0 0 18 0 0 13 3
249 91
228 91
228 147
2 1 4 0 0 0 0 10 12 0 0 2
251 147
202 147
1 4 5 0 0 0 0 8 10 0 0 2
269 171
269 166
1 3 6 0 0 0 0 9 10 0 0 2
269 135
269 140
2 0 7 0 0 0 0 12 0 0 18 2
184 147
157 147
1 1 2 0 0 0 0 11 17 0 0 4
157 202
157 204
157 204
157 197
2 0 7 0 0 0 0 17 0 0 20 2
157 161
157 147
2 5 3 0 0 0 0 16 10 0 0 4
205 62
303 62
303 153
287 153
1 2 7 0 0 0 0 16 19 0 0 4
187 62
157 62
157 147
146 147
1 1 8 0 0 0 0 19 13 0 0 2
110 147
78 147
1 2 2 0 0 0 0 15 13 0 0 3
85 202
85 157
78 157
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
402 104 439 128
412 112 428 128
2 +V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
400 179 437 203
410 187 426 203
2 -V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
34 111 61 135
39 115 55 131
2 Vi
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
432 134 469 158
442 142 458 158
2 Vo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
252 100 289 124
262 108 278 124
2 +V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
250 175 287 199
260 183 276 199
2 -V
0
9 0 0
0
0
2 V1
-0.7 -1.5 -0.02
0
0 0 0
100 0 10 10000
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2032608 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 5e-06 10
0
2163704 4421696 100 100 0 0
77 66 779 156
-4 333 798 572
545 66
779 66
779 73
779 151
0 0
0 0 0 0 0 0
12403 4
4 500 1000
1
369 149
0 3 0 0 3	0 23 0 0
6030466 4421696 100 100 0 0
77 66 767 156
-4 333 798 572
86 66
77 66
767 97
767 97
0 0
0 0 0 0 0 0
12401 0
4 20 0.5
1
324 112
0 5 0 0 3	0 23 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
