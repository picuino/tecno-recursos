CircuitMaker Text
5.6
Probes: 2
U2_6
Transient Analysis
0 677 147 65280
U2_6
AC Analysis
0 688 149 8421376
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
21 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 361
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1446 465
144179218 0
0
6 Title:
5 Name:
0
0
0
20
10 Capacitor~
219 488 153 0 2 5
0 6 4
0
0 0 848 0
6 0.01uF
-22 -18 20 -10
2 C4
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4299 0 0
2
5.89938e-315 0
0
2 +V
167 639 175 0 1 3
0 7
0
0 0 54256 180
4 -15V
3 -2 31 6
2 V6
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9672 0 0
2
5.89938e-315 5.26354e-315
0
2 +V
167 639 126 0 1 3
0 8
0
0 0 54256 0
3 15V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7876 0 0
2
5.89938e-315 5.30499e-315
0
7 Ground~
168 598 230 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6369 0 0
2
5.89938e-315 5.32571e-315
0
10 Capacitor~
219 555 153 0 2 5
0 5 4
0
0 0 848 180
6 0.01uF
-21 -18 21 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9172 0 0
2
5.89938e-315 5.34643e-315
0
8 Op-Amp5~
219 639 147 0 5 11
0 5 9 8 7 3
0
0 0 848 0
5 UA741
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 256 1 0 0 0
1 U
7100 0 0
2
5.89938e-315 5.3568e-315
0
8 Op-Amp5~
219 317 149 0 5 11
0 15 14 13 12 6
0
0 0 848 0
5 UA741
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 256 1 0 0 0
1 U
3820 0 0
2
5.89938e-315 5.36716e-315
0
10 Capacitor~
219 276 200 0 2 5
0 2 15
0
0 0 848 90
7 0.001uF
7 0 56 8
2 C1
13 -10 27 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7678 0 0
2
5.89938e-315 5.37752e-315
0
11 Signal Gen~
195 105 160 0 64 64
0 11 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162722
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V1
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 1 0 0
1 V
961 0 0
2
5.89938e-315 5.38788e-315
0
7 Ground~
168 276 232 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3178 0 0
2
5.89938e-315 5.39306e-315
0
7 Ground~
168 136 232 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3409 0 0
2
5.89938e-315 5.39824e-315
0
2 +V
167 317 128 0 1 3
0 13
0
0 0 54256 0
3 15V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3951 0 0
2
5.89938e-315 5.40342e-315
0
2 +V
167 317 177 0 1 3
0 12
0
0 0 54256 180
4 -15V
3 -2 31 6
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8885 0 0
2
5.89938e-315 5.4086e-315
0
10 Capacitor~
219 239 50 0 2 5
0 10 6
0
0 0 848 0
7 0.002uF
-25 -18 24 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3780 0 0
2
5.89938e-315 5.41378e-315
0
9 Resistor~
219 568 48 0 2 5
0 4 3
0
0 0 880 0
6 11.25k
-21 -14 21 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9265 0 0
2
5.89938e-315 5.41896e-315
0
9 Resistor~
219 648 80 0 2 5
0 9 3
0
0 0 880 0
5 22.5k
-18 -14 17 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9442 0 0
2
5.89938e-315 5.42414e-315
0
9 Resistor~
219 598 195 0 3 5
0 2 5 -1
0
0 0 880 90
5 22.5k
11 0 46 8
2 R4
22 -10 36 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9424 0 0
2
5.89938e-315 5.42933e-315
0
9 Resistor~
219 239 155 0 2 5
0 10 15
0
0 0 880 0
6 11.25k
-21 -14 21 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9968 0 0
2
5.89938e-315 5.43192e-315
0
9 Resistor~
219 326 82 0 2 5
0 14 6
0
0 0 880 0
5 22.5k
-18 -14 17 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9281 0 0
2
5.89938e-315 5.43451e-315
0
9 Resistor~
219 173 155 0 2 5
0 11 10
0
0 0 880 0
6 11.25k
-21 -14 21 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8464 0 0
2
5.89938e-315 5.4371e-315
0
23
2 0 3 0 0 4224 0 15 0 0 10 3
586 48
697 48
697 80
1 0 4 0 0 8320 0 15 0 0 6 3
550 48
517 48
517 153
1 1 2 0 0 4096 0 17 4 0 0 2
598 213
598 224
2 0 5 0 0 4096 0 17 0 0 5 2
598 177
598 153
1 1 5 0 0 4224 0 5 6 0 0 2
564 153
621 153
2 2 4 0 0 0 0 5 1 0 0 2
546 153
497 153
1 0 6 0 0 12288 0 1 0 0 18 4
479 153
458 153
458 148
375 148
1 4 7 0 0 0 0 2 6 0 0 2
639 160
639 160
1 3 8 0 0 4224 0 3 6 0 0 2
639 135
639 134
2 5 3 0 0 0 0 16 6 0 0 4
666 80
697 80
697 147
657 147
2 1 9 0 0 8320 0 6 16 0 0 4
621 141
598 141
598 80
630 80
2 0 6 0 0 4224 0 14 0 0 18 3
248 50
375 50
375 82
1 0 10 0 0 8320 0 14 0 0 15 3
230 50
206 50
206 155
1 1 11 0 0 4224 0 20 9 0 0 2
155 155
136 155
2 1 10 0 0 0 0 20 18 0 0 2
191 155
221 155
1 4 12 0 0 0 0 13 7 0 0 2
317 162
317 162
1 3 13 0 0 4224 0 12 7 0 0 2
317 137
317 136
2 5 6 0 0 0 0 19 7 0 0 4
344 82
375 82
375 149
335 149
2 1 14 0 0 8320 0 7 19 0 0 4
299 143
276 143
276 82
308 82
1 2 2 0 0 4224 0 11 9 0 0 2
136 226
136 165
1 1 2 0 0 0 0 10 8 0 0 2
276 226
276 209
2 0 15 0 0 4096 0 8 0 0 23 3
276 191
276 155
277 155
2 1 15 0 0 4224 0 18 7 0 0 4
257 155
300 155
300 155
299 155
0
0
25 0 0
0
0
2 V1
-0.7 -1.5 -0.02
0
0 0 0
50000 0 10 1e+06
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1442704 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 5e-06 10
0
1311672 4356672 100 100 0 0
77 66 777 156
-4 333 798 572
326 66
498 66
777 103
777 156
0 0
0 0 0 0 0 0
12403 1
4 500 1000
1
697 147
0 3 0 0 2	0 10 0 0
6030466 4421696 100 100 0 0
77 66 767 156
-4 333 798 572
86 66
77 66
767 97
767 97
0 0
0 0 0 0 0 0
12401 0
4 20 0.5
1
324 112
0 5 0 0 3	0 24 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
