CircuitMaker Text
5.6
Probes: 2
U1_6
Operating Point
0 361 151 65280
U1_6
AC Analysis
0 353 149 8421376
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
21 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 361
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1446 465
9961490 0
0
6 Title:
5 Name:
0
0
0
10
8 Op-Amp5~
219 317 149 0 5 11
0 5 3 8 7 3
0
0 0 80 0
5 UA741
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
4299 0 0
2
44525.4 0
0
10 Capacitor~
219 233 155 0 2 5
0 5 4
0
0 0 848 180
6 0.01uF
-22 -18 20 -10
2 C2
-8 -31 6 -23
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9672 0 0
2
44525.4 1
0
11 Signal Gen~
195 105 160 0 64 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162722
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 592 0
5 -1/1V
-18 -30 17 -22
2 Vi
-6 -31 8 -23
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 1 0 0
1 V
7876 0 0
2
44525.4 2
0
7 Ground~
168 276 232 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6369 0 0
2
44525.4 3
0
7 Ground~
168 136 232 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9172 0 0
2
44525.4 4
0
2 +V
167 317 118 0 1 3
0 8
0
0 0 53616 0
3 15V
-9 -25 12 -17
2 V1
-6 -14 8 -6
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7100 0 0
2
44525.4 5
0
2 +V
167 317 186 0 1 3
0 7
0
0 0 53616 180
4 -15V
-10 1 18 9
2 V2
-6 -1 8 7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3820 0 0
2
44525.4 6
0
10 Capacitor~
219 166 155 0 2 5
0 6 4
0
0 0 848 0
6 0.01uF
-20 -19 22 -11
2 C1
-6 -30 8 -22
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7678 0 0
2
44525.4 7
0
9 Resistor~
219 276 197 0 3 5
0 2 5 -1
0
0 0 880 90
5 22.5k
5 9 40 17
2 R1
7 -6 21 2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
961 0 0
2
44525.4 8
0
9 Resistor~
219 246 50 0 2 5
0 4 3
0
0 0 880 0
6 11.25k
-24 7 18 15
2 R2
-7 -12 7 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3178 0 0
2
44525.4 9
0
11
2 0 3 0 0 12288 0 1 0 0 2 4
299 143
277 143
277 76
375 76
2 5 3 0 0 4224 0 10 1 0 0 4
264 50
375 50
375 149
335 149
1 0 4 0 0 8320 0 10 0 0 7 3
228 50
195 50
195 155
1 1 2 0 0 4096 0 9 4 0 0 2
276 215
276 226
2 0 5 0 0 4096 0 9 0 0 6 2
276 179
276 155
1 1 5 0 0 4224 0 2 1 0 0 2
242 155
299 155
2 2 4 0 0 0 0 2 8 0 0 2
224 155
175 155
1 1 6 0 0 4224 0 8 3 0 0 2
157 155
136 155
1 4 7 0 0 4224 0 7 1 0 0 2
317 171
317 162
1 3 8 0 0 4224 0 6 1 0 0 2
317 127
317 136
1 2 2 0 0 4224 0 5 3 0 0 2
136 226
136 165
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
348 145 385 169
358 153 374 169
2 Vo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
298 90 335 114
308 98 324 114
2 +V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
329 173 366 197
339 181 355 197
2 -V
0
9 0 0
0
0
2 V1
-0.7 -1.5 -0.02
0
0 0 0
100 0 10 10000
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
5768164 1210432 100 100 0 0
0 0 0 0
0 107 161 177
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 5e-06 10
0
5309400 4421696 100 100 0 0
77 66 779 156
-4 333 798 572
545 66
311 66
779 84
779 111
0 0
0 0 0 0 0 0
12403 0
4 500 1000
1
369 149
0 3 0 0 3	0 12 0 0
6030466 4421696 100 100 0 0
77 66 767 156
-4 333 798 572
86 66
77 66
767 97
767 97
0 0
0 0 0 0 0 0
12401 0
4 20 0.5
1
324 112
0 5 0 0 3	0 12 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
