��  CCircuit��  CSerializeHack           ��  CPart�� 	 CGroupBox  D�,�             �  $ ��             �  D$ ,�             �  $ $ �                           ��� 	 CFilament��  CDummyValue  ��    1W            �?      �? W �� 	 CTerminal  ��	       �#����!@cR�e�?  �  Ti	     
   ~G����@cR�e̿    ��T           ��`   ��  ����    1W            �?      �? W �  ����        [_A�6x�
cR�e̿  �  T�i�        ������@
cR�e�?    �>T�          ��`   �� 
 CBattery9V�  �8�8    9V            "@      �? V �  �(�=        [_A�6x�cR�e�?  �  �(�=        �#����!@cR�e̿    l<��         ��   �  ��  x�x�    1W            �?      �? W �  h�}�      	 ������@cR�e̿  �  ����        |G����@cR�e�?    |>��          ��`   ��  xx    1W            �?      �? W �  h}	     
 	 ~G����@cR�e�?  �  ��	        |G����@cR�e̿    |��      #     ��`   ��  PP    1W            �?      �? W �  @U        �)#���@,�����?  �  ��        bSF���@,����п    T��(     '     ��`   ��  P�P�    1W            �?      �? W �  @�U�     	       e�]�.����п  �  ����        bSF���@.�����?    TF��     +     ��`   ��  � �     1W            �?      �? W �  � �        ؔ���!@-�����?  �  � 	        �)#���@-����п    � �� (     /     ��`   ��  � @� @    9V            "@      �? V �  � 0� E      	      e�]�.�����?  �  X 0Y E        ؔ���!@.����п    D D� �     3    ��   �  ��  8� 8�     1W            �?      �? W �  (� =�       	 xA�  @��dQ��?  �  �� ��            �Zf>��dQ�տ    <F ��      7  
   ��`   ��  �� ��     9V            "@      �? V �  �� ��            �Zf>��dQ��?  �  x� y�         ��e  "@��dQ�տ    d� �X     ;    ��   �  ��  �� ��     1W            �?      �? W �  �� ��        ��e  "@��dQ��?  �  � )�         xA�  @��dQ�տ    �F �      ?  
   ��`   ��  � � � �     1W            �?      �? W �  x � � �              "@Nð���?  �  � � �                  Nð��޿    � F � �      C  
   ��`   ��  x � x �     9V            "@      �? V �  x � y �                  Nð���?  �  P � Q �               "@Nð��޿    < � � X     G    ��   �                ���  CWire  �(�)      J�  �(��       J�  ��	      J�  ��)       J�  ���       J�  � 0A1     	 J�  @0A�      	 J�  ���       J�  A      J�  X Y 1       J�  X �       J�  �� ��        J�  x� ��       J�  x� y�        J�  �� ��       J�   � �         J�  x � �        J�  P � Q �        J�  P � y �                     �                             M    #  L      K   N         O #  # $ $ O ' S ' ( ( R + Q + , , R / U / 0 0 S 3 P 3 4 T 4 7 @ 7 8 8 V ; Y ; < X < ? W ? @ @ 7 C ] C D D Z G [ G H \ H  L K  N  M  $   3 Q P + ( , 0 ' U 4 T / 8 Y X ? W < ; V D [ G Z ] H \ C   E         �4s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 