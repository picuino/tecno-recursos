��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  '    S2      �  � �     S1      �  ����    L2      �  �a�o    L1      �  � q      L1      �  Qq a     L2      �  � Y � g     S1                    ���  CBattery��  CValue  � �%     9V         "@      �? V �� 	 CTerminal  �0 �1              "@          �  �0 �1                             �$ �<         ��      �� 	 CRailThru�  0 -1       e       "@          �  0 11              "@            , .4          ����    ��  P -Q        d                   �  P 1Q                             L .T          ����    ��  � -�       d        �          �  � 1�                             � .�          ����    ��  CSPDT��  CToggle  ��0      "   �  �                �          �  �� ��                �          �  ��	                            �� �    %      ��    ��  0-1      d                   �  011                            ,.4     )    ����    ��  -	      d        �          �  1	                            .     ,    ����    ��  � -�       d        �          �  � 1�                             � .�      /    ����    ��  � -�       d                   �  � 1�                             � .�      2    ����    !�#�  �� ��       4   �  �� �                �          �  �� ��                �          �  �� ��                             �� ��     6      ��    ��  p -q       d        �          �  p 1q                             l .t      :    ����    ��  P-Q     
 d        �          �  P1Q                            L.T     =    ����    ��  CBulb�  �P	Q     
          �          �  �P�Q               �            �D�\    A    ��      ��  p-q      d        �          �  p1q     	                       l.t     D    ����    ��  �-�      d        �          �  �1�                            �.�     G    ����    ?��  ��	�               �          �  ����               �            ����    J    ��      ��  �-�      d        �          �  �1�                            �.�     M    ����    ?��  � X � m                 �          �  � � � �                �            � l � �      P    ��      ?��  @X Am                 �          �  @� A�                �            4l L�      S    ��      ��   q 3      9V(          "@      �? V �  @ X A m               "@          �  @ � A �                �            4 l L �      W    ��      ��  CSPST#�  x 8 � X       Z   �  h 0 } 1              "@          �  � 0 � 1                �            | , � 4      \      ��                  ���  CWire  �0 1       _�  �P Q        _�  �0 �Q         _�  �0 �1        _�  �� ��       _�  �� ��        _�  �� �       _�          _�   	       _�  	      _�  �01      _�  ��1       _�  ��	      _�  �� ��       _�  �� ��        _�  �� �       _�  � �       _�  � �        _�   � �       _�  �p q       _�  �p ��        _�  �� ��       _�  PQ     
 _�  �pq      _�  �P�q       _�  �P�Q      _�  ����      _�  ����       _�  ���      _�  ��      _�  @ � A �        _�  @ � � �       _�  � 0 A1       _�  � 0 � 1       _�  � � A�       _�  � � � �        _�  @0 AY        _�  � 0 � Y        _�  @� A�        _�  @ 0 A Y        _�  @ 0 i 1                     �                              `  c  `      a      f        % % g & d & ' l ' j ) * *   i , - -   p / 0 0   o 2 3 3   6 6 r 7 u 7 8 m 8 s : ; ;   v = > >   A A v B y B w D E E   | G H H   J J } K z K } M N N   P � P Q Q � S � S T T � W � W X X ~ \ � \ ] ] �   b  c a b  e & f d e  % h g i h , k ) l j k ' n 8 m o n 2 q / r p 6 q t : s u t 7 A = x D y w x B { K z | { G J M X  ~ � � � ] � � � Q  � S � P T � � W � \            �%s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 