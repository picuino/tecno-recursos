CircuitMaker Text
5.6
Probes: 2
C2_1
Transient Analysis
0 386 187 65280
C2_1
AC Analysis
0 382 188 8421376
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 361
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
46 C:\Archivos de programa\CircuitMaker 6\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1446 465
144179218 0
0
6 Title:
5 Name:
0
0
0
12
10 Polar Cap~
219 308 35 0 2 5
0 3 6
0
0 0 848 180
6 0.01uF
-25 -18 17 -10
2 C2
-11 -28 3 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3536 0 0
2
5.89938e-315 0
0
10 Polar Cap~
219 257 181 0 2 5
0 4 6
0
0 0 848 180
6 0.01uF
-25 -18 17 -10
2 C1
-11 -28 3 -20
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4597 0 0
2
5.89938e-315 5.26354e-315
0
2 +V
167 325 249 0 1 3
0 7
0
0 0 54256 180
4 -10V
3 -2 31 6
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3835 0 0
2
44525.5 0
0
2 +V
167 325 138 0 1 3
0 8
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3670 0 0
2
44525.5 1
0
7 Ground~
168 118 275 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
44525.5 2
0
11 Signal Gen~
195 72 187 0 19 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 Vi
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9323 0 0
2
44525.5 3
0
7 Ground~
168 285 277 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
317 0 0
2
44525.5 4
0
7 Ground~
168 212 276 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3108 0 0
2
44525.5 5
0
8 Op-Amp5~
219 324 186 0 5 11
0 2 4 8 7 3
0
0 0 848 0
5 LF353
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 589827
88 0 0 256 2 1 1 0
1 U
4299 0 0
2
44525.5 6
0
9 Resistor~
219 328 86 0 2 5
0 4 3
0
0 0 880 0
3 16k
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9672 0 0
2
44525.5 7
0
9 Resistor~
219 213 231 0 3 5
0 2 6 -1
0
0 0 880 90
3 16k
12 1 33 9
2 Rr
9 -10 23 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7876 0 0
2
44525.5 8
0
9 Resistor~
219 146 182 0 2 5
0 5 6
0
0 0 880 0
2 8k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6369 0 0
2
44525.5 9
0
13
2 0 3 0 0 4096 0 10 0 0 7 2
346 86
400 86
0 1 4 0 0 4224 0 0 10 6 0 3
287 180
287 86
310 86
1 1 5 0 0 4224 0 12 6 0 0 2
128 182
103 182
2 0 6 0 0 4096 0 12 0 0 5 4
164 182
214 182
214 182
213 182
2 0 6 0 0 0 0 11 0 0 13 2
213 213
213 180
1 2 4 0 0 0 0 2 9 0 0 3
264 181
264 180
306 180
5 1 3 0 0 8320 0 9 1 0 0 4
342 186
400 186
400 35
315 35
1 4 7 0 0 4224 0 3 9 0 0 3
325 234
325 199
324 199
1 3 8 0 0 4224 0 4 9 0 0 3
325 147
325 173
324 173
1 2 2 0 0 4096 0 5 6 0 0 3
118 269
118 192
103 192
1 1 2 0 0 4224 0 7 9 0 0 3
285 271
285 192
306 192
1 1 2 0 0 0 0 8 11 0 0 4
212 270
212 255
213 255
213 249
2 2 6 0 0 8320 0 1 2 0 0 4
298 35
213 35
213 181
247 181
0
0
2073 0 1
0
0
0
0 0 0
0
0 0 0
20000 0 1 1e+06
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
4654008 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 5
0
4391674 8550464 100 100 0 0
77 66 647 246
680 74 1360 406
647 66
77 66
647 66
647 246
0 0
0 0 0 0 0 0
12401 0
4 0.001 5
1
112 179
0 9 0 0 1	0 14 0 0
1311754 4356160 100 100 0 0
77 66 647 246
680 406 1360 738
647 66
77 66
647 67
647 246
0 0
0 0 0 0 0 0
12401 0
4 30 50
1
382 186
0 11 0 0 3	0 14 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
