��  CCircuit��  CSerializeHack           ��  CPart�� 	 CGroupBox  D�,�             �  $ ��             �  D$ ,�             �  $ $ �                           ���  CBattery��  CDummyValue  0000    1.5V            �?      �? V �� 	 CTerminal  0 15        `SF����>KT�J�ؿ  �  0�1�       ؔ����h�J��?     4@�         ��   �  ��  �0�0    1.5V            �?      �? V �  � �5      
   ���  �?�_��J�ؿ  �  ����       `SF����>KT�J��?    �4��         ��   �  ��  � 0� 0    1.5V            �?      �? V �  �  � 5            `�MC>$�2R�տ  �  � �� �       tM��������dQ��?    � 4� �         ��   �  ��  �0�0    1.5V            �?      �? V �  � �5         (k�   @=KT�J�ؿ  �  ����     
  ���  �?�_��J��?    �4��         ��   �  ��  h0h0    1.5V            �?      �? V �  h i5      	   (k�   @g�J�ؿ  �  h�i�        (k�   @=KT�J��?    X4x�     "    ��   �  �� 	 CFilament�  ��    1W            �?      �? W �  ��	     	   (k�   @h�J��?  �  �		       ؔ����h�J�ؿ    ���      '  
   ��`   $��  pp    1W            �?      �? W �  `u	        F�4  @��dQ��?  �  ��	       tM��������dQ�տ    t��      +  
   ��`   ��  H 0H 0    1.5V            �?      �? V �  H  I 5         F�4  @��dQ�տ  �  H �I �        ��i  �?$�2R��?    8 4X �     /    ��   �  ��  � 0� 0    1.5V            �?      �? V �  �  � 5         ��i  �?$�2R�տ  �  � �� �          `�MC>$�2R��?    x 4� �     3    ��   �  ��  �� ��     1.5V            �?      �? V �  �� ��                �?�����п  �  �<�Q                ������?    �� �<     7    ��   �  ��  h� h�     1.5V            �?      �? V �  h� i�                @,����п  �  h<iQ              �?������?    X� x<     ;    ��   �  $��  �� ��     1W            �?      �? W �  �� ��               @,�����?  �  �� 	�                  ,����п    �> ��      ?     ��`   $��  p� p�     1W            �?      �? W �  `� u�               �?D�S�a]�?  �  �� ��                �D�S�a]ƿ    t> ��      C     ��`   ��  H � H �     1.5V            �?      �? V �  H � I �                �?D�S�a]ƿ  �  H <I Q               �D�S�a]�?    8 � X <     G    ��   �                ���  CWire   1!      J�   	�       J�  ��	�      J�  � �!     
 J�  � ��      
 J�  ����     
 J�  0�	�      J�  h�	     	 J�  � �� �      J�  �  � �       J�  �  � !      J�  � ���      J�  hi!      	 J�  	�       J�  h���      J�  � ��       J�  � �!      J�  h  � !      J�  h  i �       J�  H �i �      J�  ���       J�  H I !       J�  H a	      J�  h� ��       J�  h� i�        J�  H � a�       J�  H � I �        J�  � 	Q        J�  �P	Q       J�  hP�Q      J�  �� �Q       J�  �� ��       J�  �� �Q       J�  H P�Q                    �                             K    Q  N    M  U    V  [    P " W " # # Y ' R ' ( ( X + a + , , _ / ` / 0 0 ^ 3 \ 3 4 4 S 7 j 7 8 8 g ; c ; < < h ? b ? @ @ f C d C D D k G e G H H l L  K M  L O  N P  O  X W ' 4 T U S T   _ R " ( Q # Z [ Y Z  ] 3 \ ^ 0 ] , V a / ` + c ? b ; e C d G @ g 8 f < i j h i 7 D l H k   5         �4s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 