��  CCircuit��  CSerializeHack           ��  CPart�� 	 CGroupBox  $ P�             �  $  D             �  D ,D             �  DT,,                           ��� 	 CFilament��  CDummyValue  HH    1W            �?      �? W �� 	 CTerminal  8M	     	           Nð��޿  �  ��	             "@Nð���?    L��        
   ��`   ��  H�H�    1W            �?      �? W �  8�M�     	           Nð��޿  �  ����             "@Nð���?    LF��       
   ��`   ��  H(H(    1W            �?      �? W �  8(M)     	           Nð��޿  �  �(�)             "@Nð���?    L��@       
   ��`   ��  H�H�    1W            �?      �? W �  8�M�     	           Nð��޿  �  ����             "@Nð���?    Lf��       
   ��`   �� 
 CBattery9V�  ����    9V            "@      �? V �  ����      	          Nð���?  �  x�y�              "@Nð����    d��x     #    ��   �  ��   � �    1W            �?      �? W �  �%�               �Nð��޿  �  ����             "@Nð���?    $V��     '  
   ��`   ��   0 0    1W            �?      �? W �  0%1               �Nð��޿  �  �0�1             "@Nð���?    $��H     +  
   ��`    ��  x �x �    9V            "@      �? V �  x �y �               ��U�D��?  �  P �Q �              "@�U�D���    < �� x     /    ��   �  ��   � �    1W            �?      �? W �  �%�               �Nð��޿  �  ����             "@Nð���?    $n��     3  
   ��`   ��   �  �     1W            �?      �? W �  � %�                  Nð��޿  �  �� ��              "@Nð���?    $. ��      7  
   ��`    ��  x � x �     9V            "@      �? V �  x � y �                  Nð���?  �  P � Q �               "@Nð��޿    < � � 8     ;    ��   �  ��  H� H�     1W            �?      �? W �  8� M�             e�]�Nð��޿  �  �� ��        ؔ���!@Nð���?    L. ��      ?  
   ��`    ��  �� ��     9V            "@      �? V �  �� ��             e�]�Nð���?  �  x� y�         ؔ���!@Nð���    d� �8     C    ��   �  ��  H� H�     1W            �?      �? W �  8� M�             e�]�Nð��޿  �  �� ��        ؔ���!@Nð���?    L� �     G  
   ��`                 ���  CWire  �(��       J�  ���	       J�  ����      	 J�  ��9�     	 J�  8�9)      	 J�  8(9�      	 J�  8�9	      	 J�  ���)       J�  �`��       J�  x`�a      J�  x`y�       J�  �0��       J�  0�       J�  �1       J�  P `Q �       J�  P `�a      J�  x �y �       J�  x ��      J�  ���1       J�  �`��       J�  x � �        J�  x � y �         J�  �  ��        J�  P   �!       J�  P   Q �        J�  �� 9�       J�  �� ��        J�  �  ��        J�  x  �!       J�  x  y�        J�  8� 9�        J�  �� ��                      �                             Q    L  Q    L  O    R  O    R # M # $ U $ ' W ' ( ( V + W + , , ] / [ / 0 Y 0 3 \ 3 4 4 ] 7 _ 7 8 8 a ; ` ; < c < ? d ? @ @ f C e C D h D G i G H H j   K  N # M  N P   P  S K T  U S T $ , ( X ' 3 + Z 0 Y ^ \ / [ X ^ V Z 4 ` 7 _ ; b 8 c a b < e i d C g j h f g D ? G @ H  
 9        �4s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 