��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  �Y	g    L1      �  ��	�    L2      �  � *�     S1      �  *    S2      �  � A � O     S1      �  � � � �     L1      �  A� Q�     L2      �  YA jO     S2                    ��� 	 CRailThru�� 	 CTerminal  0�E�      d                   �  4�I�               �            2�F�         ����    ��  CBulb�  �!�                          �  ����               �            �|�        ��      ��  0�E�      d        �          �  4�I�                            2�F�         ����    ��  0hEi      d        �          �  4hIi                            2dFl         ����    ��  H!I               �          �  �H�I               �            �<T    !    ��      ��  0HEI      d        �          �  4HII                            2DFL     $    ����    ��  0h Ei       d        �          �  4h Ii                             2d Fl      '    ����    ��  CSPDT��  CToggle  �� �       *   �  � �                �          �  �� ��                �          �  �� ��                             �| �     -      ��    ��  0� E�       d                   �  4� I�                             2� F�      1    ����    ��  0� E�       d        �          �  4� I�                             2� F�      4    ����    ��  0 E      d        �          �  4 I                            2� F     7    ����    ��  0(E)      d                   �  4(I)                            2$F,     :    ����    )�+�  �(      <   �  � �                �          �  �� ��      	          �          �  � �                            ��     >      ��    ��  0� E�      	 d        �          �  4� I�      
                       2� F�      B    ����    ��  0H EI        d                   �  4H II                             2D FL      E    ����    ��  0( E)       e       "@          �  4( I)              "@            2$ F,      H    ����    ��  CBattery��  CValue  �      9V         "@      �? V �  �( )              "@          �  �( �)                             � �4     N    ��      ��  CSPST+�  � 8 � X       Q   �  � T � i                �          �  � ( � =               "@            � < � T     S      ��    ��  � h � }        	        �          �  � � � �                             � | � �      V    ��      ��  0h 1}        	        �          �  0� 1�                             $| <�      Y    ��      P�+�  88 XX       [   �  0T 1i                �          �  0( 1=               "@            ,< 4T     ]      ��    J�L�   Q 3 _     9V(          "@      �? V �  @ 8 A M               "@          �  @ d A y                             4 L L d      a    ��                    ���  CWire   �1�      d�  ��1�      d�  ����       d�  ����      d�  �H�I      d�  �H�i       d�  �h1i      d�   H1I      d�  �� ��       d�  �h ��        d�  �h 1i       d�  � )�       d�  (� )�        d�  (� 1�       d�  �� 1�       d�  �� ��        d�  �� ��       d�  � �      d�  � �)       d�  �(1)      d�  ( 1      d�  (� )       d�  � )�       d�  �� 1�      	 d�  �� ��       	 d�  �� ��      	 d�  �( �)        d�  �( �I         d�  �H 1I        d�  ( 1)       d�  � � 1�       d�  @ � � �       d�  @ x A �        d�  � ( 1)       d�  @ ( � )       d�  @ ( A 9                      �                            e        e  h  f      k      ! ! l " i " l $ % %   o ' ( (   - - p . m . / u / s 1 2 2   r 4 5 5   y 7 8 8   x : ; ;   > > { ? ~ ? @ v @ | B C C   � E F F   � H I I   N N � O  O S S V T � T V S V W W � Y ] Y Z Z � ] ] Y ^ � ^ a � a b b �   g  h f g  j " i k j  ! $ n . o m n ' - q p r q 4 t 1 u s t / w @ v x w : z 7 { y > z } B | ~ } ? � O  � � E N H W Z � � b � T ^ � � � a   K         �%s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 