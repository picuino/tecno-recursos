��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  ya�o    L1      �  y���    L2      �  �� ��     S1      �  ��'    S2      �  � Y � g     L1      �  � Y � g     S1                    ��� 	 CRailThru�� 	 CTerminal  ����      d                   �  ����               �            ����         ����    ��  CBulb�  ����                          �  `�u�               �            t���        ��      ��  ����      d        �          �  ����                            ����         ����    ��  �p�q      d        �          �  �p�q                            �l�t         ����    ��  �P�Q               �          �  `PuQ               �            tD�\        ��      ��  �P�Q      d        �          �  �P�Q                            �L�T     "    ����    ��  �p �q       d        �          �  �p �q                             �l �t      %    ����    ��  CSPDT��  CToggle  h� ��       (   �  �� ��                �          �  X� m�                �          �  X� m�                             l� ��     +      ��    ��  �� ��       d                   �  �� ��                             �� ��      /    ����    ��  �� ��       d        �          �  �� ��                             �� ��      2    ����    ��  ��	     
 d        �          �  ��	                            ��     5    ����    ��  �0�1      d                   �  �0�1                            �,�4     8    ����    '�)�  h�0      :   �  � �     
          �          �  X� m�                �          �  Xm	                            l� �    <      ��    ��  �� ��       d        �          �  �� ��      	                       �� ��      @    ����    ��  �P �Q        d                   �  �P �Q                             �L �T      C    ����    ��  �0 �1       e       "@          �  �0 �1              "@            �, �4      F    ����    ��  CBattery��  CValue  \ �%     9V         "@      �? V �  |0 �1              "@          �  P0 e1                             d$ |<     L    ��      H�J�   Y 3 g     9V(          "@      �? V �  @ @ A U               "@          �  @ l A �                �            4 T L l      P    ��      ��  CSPST)�  x 0 � P       S   �  h ( } )              "@          �  � ( � )                �            | $ � ,      U      ��    ��  � @ � U                 �          �  � l � �                �            � T � l      X    ��                    ���  CWire  ����      [�  @���      [�  @�A�       [�  @�a�      [�  @PaQ      [�  @PAq       [�  @p�q      [�  �P�Q      [�  @� Y�       [�  @p A�        [�  @p �q       [�  �� ��       [�  �� ��        [�  �� ��       [�  @� ��       [�  @� A�        [�  @� Y�       [�  @Y	      [�  @A1       [�  @0�1      [�  ��	     
 [�  � �	      
 [�  � �     
 [�  @� ��       [�  @� A�        [�  @� Y�       [�  @0 Q1        [�  @0 AQ         [�  @P �Q        [�  �0 �1       [�  @ ( i )       [�  @ ( A A        [�  � ( � )       [�  � ( � A        [�  @ � A �        [�  @ � � �       [�  � � � �                      �                            \        \  _  ]      b        c   `   c " # #   f % & &   + + g , d , - l - j / 0 0   i 2 3 3   p 5 6 6   o 8 9 9   < < r = u = > m > s @ A A   x C D D   y F G G   L L y M v M P { P Q Q ~ U z U V V | X } X Y Y �   ^  _ ] ^  a   ` b a   " e , f d e % + h g i h 2 k / l j k - n > m o n 8 q 5 r p < q t @ s u t = w M v x w C L F { U z P V } | X Q  ~ � Y    I         �%s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 