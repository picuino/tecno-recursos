CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1446 465
9961490 0
0
6 Title:
5 Name:
0
0
0
9
2 +V
167 190 121 0 1 3
0 6
0
0 0 53856 0
2 5V
-8 -22 6 -14
3 Vi2
-9 -13 12 -5
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6343 0 0
2
5.89977e-315 5.26354e-315
0
2 +V
167 190 64 0 1 3
0 7
0
0 0 53856 0
2 5V
-8 -22 6 -14
3 Vi1
-10 -13 11 -5
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7376 0 0
2
5.89977e-315 5.30499e-315
0
2 +V
167 292 111 0 1 3
0 8
0
0 0 53344 0
3 15V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9156 0 0
2
5.89977e-315 5.32571e-315
0
2 +V
167 292 186 0 1 3
0 9
0
0 0 53344 180
4 -15V
-12 12 16 20
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5776 0 0
2
5.89977e-315 5.34643e-315
0
7 Ground~
168 262 191 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7207 0 0
2
5.89977e-315 5.3568e-315
0
8 Op-Amp5~
219 292 144 0 5 11
0 2 4 8 9 3
0
0 0 64 0
5 LF353
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 589828
88 0 0 256 2 1 1 0
1 U
4459 0 0
2
5.89977e-315 5.36716e-315
0
9 Resistor~
219 224 80 0 3 5
0 7 4 1
0
0 0 608 0
2 1k
-7 -14 7 -6
2 R1
-6 -14 8 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3760 0 0
2
5.89977e-315 5.38788e-315
0
9 Resistor~
219 308 80 0 2 5
0 4 3
0
0 0 608 0
2 2k
-7 -14 7 -6
2 RF
-6 -14 8 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
754 0 0
2
5.89977e-315 5.39306e-315
0
9 Resistor~
219 225 138 0 3 5
0 6 4 1
0
0 0 608 0
2 1k
-7 -14 7 -6
2 R2
-7 -13 7 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9767 0 0
2
5.89977e-315 5.39824e-315
0
10
0 0 0 0 0 0 0 0 0 10 7 2
262 138
262 80
0 0 3 0 0 4096 0 0 0 9 0 2
341 144
375 144
1 1 6 0 0 4224 0 1 9 0 0 3
190 130
190 138
207 138
1 1 2 0 0 8320 0 6 5 0 0 3
274 150
262 150
262 185
1 1 7 0 0 4224 0 2 7 0 0 3
190 73
190 80
206 80
1 3 8 0 0 4224 0 3 6 0 0 2
292 120
292 131
2 1 4 0 0 16 0 7 8 0 0 2
242 80
290 80
1 4 9 0 0 4224 0 4 6 0 0 2
292 171
292 157
2 5 3 0 0 8320 0 8 6 0 0 4
326 80
341 80
341 144
310 144
2 2 4 0 0 0 0 9 6 0 0 2
243 138
274 138
3
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
358 127 379 145
362 131 374 143
2 Vo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
282 86 307 110
286 90 302 106
2 +V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
283 182 308 206
287 186 303 202
2 -V
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
100 1 0.1 1e+06
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2032918 1210432 100 100 0 0
0 0 0 0
486 365 647 435
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 10
1
334 144
0 2 0 0 3	0 9 0 0
2098462 8550464 100 100 0 0
77 66 377 156
400 74 800 322
377 66
77 66
377 66
377 156
0 0
0 0 0 0 0 0
12401 0
4 0.001 10
1
340 144
0 2 0 0 1	0 11 0 0
3540064 4356160 100 100 0 0
77 66 371 156
400 322 799 570
371 66
77 66
371 66
371 156
0 0
0 0 0 0 0 0
12403 0
4 0.3 5
1
334 144
0 2 0 0 3	0 9 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
