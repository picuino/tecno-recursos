��  CCircuit��  CSerializeHack           ��  CPart  0   0       ���  CBattery��  CValue   � ; �     9V(          "@      �? V �� 	 CTerminal  H � I �               "@          �  H � I �                             < � T �          ��      ��  CBulb�  � � � �                 �          �  � � � �                              � � � �          ��      ��  CSPST��  CToggle  � ( � H          �  p   � !              "@          �  �   � !                �            �  � $            ��    ��  � 0 � E                 �          �  � \ � q                             � D � \          ��      �
�   I ; W     9V(          "@      �? V �  H 0 I E               "@          �  H \ I q                            < D T \          ��      �� 	 CPushMake��  CKey  � � � �       !   �  p � � �              "@          �  � � � �                �            � � � �      $      ��    ��  �  � 5              "@
ףp=
�?  �  � L� a                
ףp=
��    � 4� L     '  
 ��      �
�   9; G    9V(          "@      �? V �  H  I 5              "@
ףp=
��  �  H LI a               
ףp=
�?    < 4T L     +    ��      �� 
 CPushBreak"�  � � 6      .   �  p �              "@
ףp=
�?  �  � �              "@
ףp=
��    � �      0      ��      0   0       ���  CWire  H � � �        3�  �   � !       3�  �   � 1        3�  H p � q       3�  H   I 1        3�  H   q !       3�  � � � �       3�  � � � �        3�  H � q �       3�  H � I �        3�  H `� a      3�  � �       3�  � � !       3�  H q       3�  H I !         0   0       �  0   0         0   0        =    4  ;    4  9    5  6    7  8    7 $ < $ % % : ' @ ' ( ( > + B + , , > 0 A 0 1 1 ?    6 5    9  8  % ; :  = $ <  , ( 1 @ ? ' B 0 A +  	 	         �5s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 