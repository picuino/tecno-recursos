��  CCircuit��  CSerializeHack           ��  CPart              ��� 
 CCapacitor��  CValue  ����    1�F   ���ư>      �?�F �� 	 CTerminal  ����        y����!��M���\l�>  �  ����        %(Or��w?^ ��Vl��    ����       ��      U
+j����
�  D�l�    1�F   ���ư>      �?�F �  d�y�       >�v���\"\l��  �  8�M�      	 �m�q��-�����>    L�d�       ��      - 3%�$Ѿ�
�  �,�    1�F   ���ư>      �?�F �  $�9�       �m�q����3b���  �  ���      	 y����!��8���@�>    �$�       ��      �dT)+�����  CVSlide��  CSlider  IDXl    
�   QH_    0V(          $@         V    �  dXyY                z���\r�=    \Td\         ����     �� 	 CResistor
�  �F�T    10M       �cA      �?M  �  �X�Y     
   ��l�%2?z���\r�=  �  xX�Y      	         z���\r��    �T�\         ��      ��  C741��  COpampSupply�� 
 CDummyPart  D0R    &�  o0}      XX    9V            "@      �? V       "�      �? V # �  �XY     
   ��l�%2?          �  �hi                          �  $`9a       >�v��� ��-��>    R$o     )      ��    �
�  ($    10M       �cA      �?M  �  $(9)       >�v���n8Ǟl��  �  �()     
   ��l�%2?n8Ǟl�>    $$,    .    ��      �
�  ����    100k          j�@      �?k  �  ����       	 y����!��L�P�N���  �  ����     	           L�P�N��>    ����     2    ��      �
�  �3�    100k          j�@      �?k  �  8�9�       	 �m�q��3����j�  �  8�9�                3����j�>    4�<�     6    ��      ��  CEarth�  ����      	 	         L�P�N���    ���     :    ��      8��  8�9�       	         3����j�    +�C�     <    ��      �
�  �y��    10k          ��@      �?k  �  �`�u      
   ��l�%2?_ ��Vl��  �  ����      	 %(Or��w?_ ��Vl�>    �t��     ?    ��      8��  �h�}       	                     �|�     B    ��                    ���  CWire  @(Aa       D�  �X�a      
 D�  �(�)     
 D�  �(�Y      
 D�  �X�Y     
 D�  8(A)      D�  8`Aa      D�  @`�a      D�  �`��       D�  x���      D�  �X�Y     
               ���  CProbe  �Q�`       L                                      2  @    N  6          !     F !  ! % % ) I ) * B * + + K . . J / G / 2  2 3 3 : 6  6 7 7 < : 3 : < 7 < ? F ? @ @  B * B J L O ? H / G I O ) . E + E K M L N  M   H           �%s�        @     +        @            @    "V  (      �                
          @      �? V        �      �? V         
         $@      �? V               �? V                 @      �? s 