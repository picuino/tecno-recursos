CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1446 465
9961490 0
0
6 Title:
5 Name:
0
0
0
7
10 Op-Amp5:A~
219 293 144 0 5 11
0 7 4 6 5 3
0
0 0 64 0
5 LF353
19 -25 54 -17
2 U1
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 122
88 0 0 0 2 1 1 0
1 U
9968 0 0
2
44500.6 0
0
2 +V
167 293 184 0 1 3
0 5
0
0 0 53344 180
3 -1V
-11 2 10 10
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9281 0 0
2
44500.6 1
0
2 +V
167 293 108 0 1 3
0 6
0
0 0 53344 0
3 15V
-10 -22 11 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8464 0 0
2
44500.6 2
0
7 Ground~
168 248 255 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7168 0 0
2
44500.6 3
0
2 +V
167 193 118 0 1 3
0 7
0
0 0 53856 0
4 -.2V
-14 -22 14 -14
2 Vi
-6 -14 8 -6
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3171 0 0
2
44500.6 4
0
9 Resistor~
219 292 203 0 2 5
0 4 3
0
0 0 608 0
2 1k
-7 -14 7 -6
2 RF
-6 6 8 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 12147832
82 0 0 0 1 0 0 0
1 R
4139 0 0
2
44500.6 5
0
9 Resistor~
219 248 227 0 3 5
0 2 4 -1
0
0 0 608 90
2 1k
8 0 22 8
2 R1
6 -4 20 4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 26
82 0 0 0 1 0 0 0
1 R
6435 0 0
2
44500.6 6
0
8
2 0 3 0 0 8320 0 6 0 0 5 3
310 203
331 203
331 144
1 0 4 0 0 4112 0 6 0 0 3 2
274 203
248 203
2 2 4 0 0 8320 0 1 7 0 0 3
275 150
248 150
248 209
1 1 2 0 0 4224 0 7 4 0 0 4
248 245
248 254
248 254
248 249
5 0 3 0 0 0 0 1 0 0 0 2
311 144
363 144
1 4 5 0 0 4224 0 2 1 0 0 2
293 169
293 157
1 3 6 0 0 4224 0 3 1 0 0 2
293 117
293 131
1 1 7 0 0 8320 0 5 1 0 0 3
193 127
193 138
275 138
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
282 84 307 108
286 88 302 104
2 +V
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
345 126 366 144
349 130 361 142
2 Vo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
281 178 308 202
286 182 302 198
2 -V
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1705266 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 10
1
335 144
0 2 0 0 3	0 9 0 0
1967280 8550464 100 100 0 0
77 66 767 156
0 322 800 570
767 66
77 66
767 66
767 156
0 0
0 0 0 0 0 0
12385 0
4 1e-06 10
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
