��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  � Y � g     S1      �  � Y � g     S2      �  Yq i     L1      �  �a	o    L1      �  ��	�    L2      �  � *�     S1      �  *'    S2                    ���  CSPST��  CToggle  x 8 � X          �� 	 CTerminal  h 0 } 1              "@          �  � 0 � 1                �            | , � 4            ��    ��  � 8  X          �  � 0 � 1                �          �  � 0 1                �            � , � 4            ��    ��  CBulb�  HX Im                 �          �  H� I�                              <l T�          ��      ��  CBattery��  CValue   q 3      9V(          "@      �? V �  @ X A m               "@          �  @ � A �                             4 l L �      #    ��      �� 	 CRailThru�  0�E�      d        �          �  4�I�                            2�F�     '    ����    ��  �!�               �          �  ����               �            ���    *    ��      %��  0�E�      d        �          �  4�I�                            2�F�     -    ����    %��  0pEq      d        �          �  4pIq                            2lFt     0    ����    ��  P!Q               �          �  �P�Q               �            �D\    3    ��      %��  0PEQ      d        �          �  4PIQ                            2LFT     6    ����    %��  0p Eq       d        �          �  4p Iq                             2l Ft      9    ����    ��  CSPDT�  �� �       <   �  � �                �          �  �� ��                �          �  �� ��                             �� �     >      ��    %��  0� E�       d                   �  4� I�                             2� F�      B    ����    %��  0� E�       d        �          �  4� I�                             2� F�      E    ����    %��  0E	      d        �          �  4I	     
                       2F     H    ����    %��  00E1      d                   �  40I1     	                       2,F4     K    ����    ;��  �0      M   �                  �          �  �� ��                �          �  ��	                            ��     O      ��    %��  0� E�       d        �          �  4� I�                             2� F�      S    ����    %��  0P EQ       d                   �  4P IQ                             2L FT      V    ����    %��  00 E1       e       "@          �  40 I1              "@            2, F4      Y    ����    �!�  � %     9V         "@      �? V �  �0 1              "@          �  �0 �1                            �$ �<     ]    ��                    ���  CWire  H0 IY        `�  0 I1       `�  � 0 � 1       `�  @ 0 i 1       `�  @ 0 A Y        `�  H� I�         `�  @ � I�        `�  @ � A �         `�   �1�      `�  ��1�      `�  ����       `�  ����      `�  �P�Q      `�  �P�q       `�  �p1q      `�   P1Q      `�  �� ��       `�  �p ��        `�  �p 1q       `�  � )�       `�  (� )�        `�  (� 1�       `�  �� 1�       `�  �� ��        `�  �� ��       `�  ��	      `�  ��1       `�  �011      `�  (1	      `�  ( )	       `�   )      `�  �� 1�       `�  �� ��        `�  �� ��       `�  �0 �1       `�  �0 �Q        `�  �P 1Q       `�  0 11                     �                             d    c  c    b  a    f # e # $ $ h i ' ( (   * * i + l + j - . .   o 0 1 1   3 3 p 4 m 4 p 6 7 7   s 9 : :   > > t ? q ? @ y @ w B C C   v E F F   } H I I   | K L L   O O  P � P Q z Q � S T T   � V W W   � Y Z Z   ] ] � ^ � ^ b   a   e  d #  g h f $ g * ' k - l j k + n 4 m o n 0 3 6 r ? s q r 9 > u t v u E x B y w x @ { Q z | { K ~ H  } O ~ � S � � � P � ^ � � � V ] Y             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 