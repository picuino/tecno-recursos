CircuitMaker Text
5.6
Probes: 2
Vo
Transient Analysis
0 278 116 8421376
Vi_1
Transient Analysis
1 113 109 4227327
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 361
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1446 465
9961490 0
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 201 180 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3656 0 0
2
5.90006e-315 0
0
10 Capacitor~
219 176 108 0 2 5
0 6 4
0
0 0 832 0
6 0.01uF
-22 -18 20 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3131 0 0
2
5.90006e-315 5.26354e-315
0
11 Terminal:A~
194 290 114 0 1 3
0 3
0
0 0 57568 180
2 Vo
-7 -13 7 -5
2 J1
-7 -23 7 -15
0
3 Vo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
6772 0 0
2
5.90006e-315 5.30499e-315
0
2 +V
167 243 76 0 1 3
0 8
0
0 0 53600 0
3 15V
-10 -14 11 -6
3 Vi4
-10 -24 11 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9557 0 0
2
5.90006e-315 5.32571e-315
0
2 +V
167 243 160 0 1 3
0 9
0
0 0 53600 180
4 -15V
-14 -1 14 7
3 Vi3
-10 0 11 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5789 0 0
2
5.90006e-315 5.34643e-315
0
7 Ground~
168 111 180 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7328 0 0
2
5.90006e-315 5.3568e-315
0
8 Op-Amp5~
219 243 114 0 5 11
0 5 4 8 9 3
0
0 0 64 0
5 LF353
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 589828
88 0 0 0 2 1 1 0
1 U
4799 0 0
2
5.90006e-315 5.36716e-315
0
11 Signal Gen~
195 75 113 0 33 64
0 7 2 5 86 -8 8 9 0 0
0 0 0 0 0 0 0 1016028201 0 0
992204554 1045220557 1000593162 0 1005961871 -1102263091 1008981770 0 1011666125 1045220557
1014350479 0 1016028201 -1102263091
20
0 0.0175 0 0 0.0025 0.2 0.005 0 0.0075 -0.2
0.01 0 0.0125 0.2 0.015 0 0.0175 -0.2 0 0
0
0 0 832 0
11 -200m/200mV
-39 -31 38 -23
2 Vi
-7 -40 7 -32
0
0
84 %D %1 %2 DC 0 PWL( 0 0 2.5m 200m 5m 0 7.5m -200m 10m 0 12.5m 200m 15m 0 17.5m -200m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9196 0 0
2
5.90006e-315 5.37752e-315
0
9 Resistor~
219 244 35 0 2 5
0 4 3
0
0 0 864 0
4 100k
-13 -14 15 -6
2 Rf
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3857 0 0
2
5.90006e-315 5.38788e-315
0
9 Resistor~
219 201 148 0 3 5
0 2 5 -1
0
0 0 864 90
2 5k
-23 -1 -9 7
2 R2
-21 -12 -7 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7125 0 0
2
5.90006e-315 5.39306e-315
0
9 Resistor~
219 134 108 0 2 5
0 7 6
0
0 0 864 0
3 10k
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3641 0 0
2
5.90006e-315 5.39824e-315
0
11
2 1 3 0 0 8320 0 9 3 0 0 3
262 35
284 35
284 114
1 0 4 0 0 8320 0 9 0 0 5 3
226 35
201 35
201 108
1 1 2 0 0 4096 0 10 1 0 0 2
201 166
201 174
1 2 5 0 0 4224 0 7 10 0 0 3
225 120
201 120
201 130
2 2 4 0 0 0 0 2 7 0 0 2
185 108
225 108
1 2 6 0 0 4224 0 2 11 0 0 2
167 108
152 108
1 1 7 0 0 4224 0 11 8 0 0 2
116 108
106 108
5 1 3 0 0 0 0 7 3 0 0 2
261 114
284 114
3 1 8 0 0 4224 0 7 4 0 0 2
243 101
243 85
1 4 9 0 0 4224 0 5 7 0 0 2
243 145
243 127
2 1 2 0 0 8320 0 8 6 0 0 3
106 118
111 118
111 174
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.0175 7e-05 7e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2425688 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 10
0
2491180 8550464 100 100 0 0
77 66 767 156
0 322 800 570
472 66
77 66
767 66
767 156
0 0
0 0 0 0 0 0
12401 0
4 0.01 10
2
116 108
0 7 0 0 1	0 7 0 0
272 114
0 3 0 0 1	0 8 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
