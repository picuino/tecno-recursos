CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
7
10 Polar Cap~
219 243 44 0 2 5
0 4 3
0
0 0 576 0
3 1uF
-9 -18 12 -10
1 C
-5 -19 2 -11
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5130 0 0
2
5.89977e-315 0
0
2 +V
167 135 90 0 1 3
0 5
0
0 0 53856 0
3 10V
-11 -22 10 -14
2 Vi
-7 -15 7 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
5.89977e-315 5.26354e-315
0
7 Ground~
168 200 156 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3124 0 0
2
5.89977e-315 5.30499e-315
0
2 +V
167 243 76 0 1 3
0 6
0
0 0 53344 0
3 15V
-10 -14 11 -6
3 Vi4
-10 -24 11 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3421 0 0
2
5.89977e-315 5.32571e-315
0
2 +V
167 243 160 0 1 3
0 7
0
0 0 53344 180
4 -15V
-14 -1 14 7
3 Vi3
-10 0 11 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
5.89977e-315 5.34643e-315
0
8 Op-Amp5~
219 243 114 0 5 11
0 2 4 6 7 3
0
0 0 64 0
5 LF353
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 589828
88 0 0 0 2 1 1 0
1 U
5572 0 0
2
5.89977e-315 5.3568e-315
0
9 Resistor~
219 167 108 0 3 5
0 5 4 1
0
0 0 608 0
4 100k
-13 -14 15 -6
1 R
-3 -12 4 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8901 0 0
2
5.89977e-315 5.36716e-315
0
8
0 0 3 0 0 4096 0 0 0 6 0 2
283 114
315 114
1 0 4 0 0 8320 0 1 0 0 4 3
232 44
201 44
201 108
1 1 5 0 0 4224 0 7 2 0 0 3
149 108
135 108
135 99
2 2 4 0 0 0 0 7 6 0 0 2
185 108
225 108
1 1 2 0 0 8320 0 6 3 0 0 3
225 120
200 120
200 150
5 2 3 0 0 8320 0 6 1 0 0 4
261 114
283 114
283 44
249 44
3 1 6 0 0 4224 0 6 4 0 0 2
243 101
243 85
1 4 7 0 0 4224 0 5 6 0 0 2
243 145
243 127
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
229 55 256 79
234 59 250 75
2 +V
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
296 95 317 113
300 99 312 111
2 Vo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
230 152 255 176
234 156 250 172
2 -V
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.0175 7e-05 7e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2425688 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 10
0
2491180 8550464 100 100 0 0
77 66 767 156
0 322 800 570
472 66
77 66
767 66
767 156
0 0
0 0 0 0 0 0
12401 0
4 0.01 10
2
116 108
0 7 0 0 1	0 9 0 0
272 114
0 3 0 0 1	0 6 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
