��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  � �     L2      �  I W     L1      �  � Y � g     S1      �  �a�o    L1      �  ����    L2      �  �� ��     S1      �  ��'    S2                    ���  CBulb�� 	 CTerminal  � p � �        	        �          �  � � � �                              � � � �          ��      ��  � 0 � E                 �          �  � \ � q                �            � D � \          ��      ��  CSPST��  CToggle  x 8 � X          �  h 0 } 1              "@          �  � 0 � 1                �            | , � 4            ��    ��  CBattery��  CValue   q 3      9V(          "@      �? V �  @ X A m               "@          �  @ � A �                             4 l L �      "    ��      �� 	 CRailThru�  ����      d        �          �  ����                            ����     &    ����    ��  ����               �          �  ����               �            ����    )    ��      $��  ����      d        �          �  ����                            ����     ,    ����    $��  �p�q      d        �          �  �p�q                            �l�t     /    ����    ��  �P�Q               �          �  �P�Q               �            �D�\    2    ��      $��  �P�Q      d        �          �  �P�Q                            �L�T     5    ����    $��  �p �q       d        �          �  �p �q                             �l �t      8    ����    ��  CSPDT�  �� ��       ;   �  �� ��                �          �  x� ��                �          �  x� ��                             �� ��     =      ��    $��  �� ��       d                   �  �� ��                             �� ��      A    ����    $��  �� ��       d        �          �  �� ��                             �� ��      D    ����    $��  ��	      d        �          �  ��	     
                       ��     G    ����    $��  �0�1      d                   �  �0�1     	                       �,�4     J    ����    :��  ��0      L   �  � �               �          �  x� ��                �          �  x�	                            �� �    N      ��    $��  �� ��       d        �          �  �� ��                             �� ��      R    ����    $��  �P �Q       d                   �  �P �Q                             �L �T      U    ����    $��  �0 �1       e       "@          �  �0 �1              "@            �, �4      X    ����    � �  | �%     9V         "@      �? V �  �0 �1              "@          �  p0 �1                            �$ �<     \    ��                    ���  CWire  @ � � �        _�  @ � A �         _�  � 0 � 1       _�  @ 0 i 1       _�  @ 0 A Y        _�  ����      _�  `���      _�  `�a�       _�  `���      _�  `P�Q      _�  `Paq       _�  `p�q      _�  �P�Q      _�  `� y�       _�  `p a�        _�  `p �q       _�  �� ��       _�  �� ��        _�  �� ��       _�  `� ��       _�  `� a�        _�  `� y�       _�  `y	      _�  `a1       _�  `0�1      _�  ��	      _�  � �	       _�  � �      _�  `� ��       _�  `� a�        _�  `� y�       _�  `0 q1       _�  `0 aQ        _�  `P �Q       _�  �0 �1                     �                                 `  b      c    b " d " # # a e & ' '   ) ) e * h * f , - -   k / 0 0   2 2 l 3 i 3 l 5 6 6   o 8 9 9   = = p > m > ? u ? s A B B   r D E E   y G H H   x J K K   N N { O ~ O P v P | R S S   � U V V   � X Y Y   \ \ � ]  ] a  # `   d  c " ) & g , h f g * j 3 i k j / 2 5 n > o m n 8 = q p r q D t A u s t ? w P v x w J z G { y N z } R | ~ } O � ]  � � U \ X            �%s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 