CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
10
2 +V
167 178 134 0 1 3
0 8
0
0 0 53856 0
2 1V
-8 -22 6 -14
3 Vi1
-8 -13 13 -5
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5130 0 0
2
44500.7 0
0
7 Ground~
168 254 205 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
391 0 0
2
44500.7 1
0
2 +V
167 178 58 0 1 3
0 5
0
0 0 53856 0
2 1V
-8 -22 6 -14
3 Vi2
-9 -12 12 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
44500.7 2
0
2 +V
167 292 116 0 1 3
0 6
0
0 0 53344 0
3 15V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3421 0 0
2
44500.7 3
0
2 +V
167 292 182 0 1 3
0 9
0
0 0 53344 180
4 -15V
-12 12 16 20
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
44500.7 4
0
8 Op-Amp5~
219 292 144 0 5 11
0 4 7 6 9 3
0
0 0 64 0
5 LF353
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 589828
88 0 0 0 2 1 1 0
1 U
5572 0 0
2
44500.7 5
0
9 Resistor~
219 254 176 0 3 5
0 2 4 -1
0
0 0 608 90
2 1k
8 0 22 8
2 R2
-17 -5 -3 3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8901 0 0
2
44500.7 6
0
9 Resistor~
219 218 75 0 3 5
0 5 7 1
0
0 0 608 0
2 1k
-7 -14 7 -6
2 R3
-7 -14 7 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7361 0 0
2
44500.7 7
0
9 Resistor~
219 298 75 0 2 5
0 7 3
0
0 0 608 0
2 1k
-7 -14 7 -6
2 RF
-7 -13 7 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4747 0 0
2
44500.7 8
0
9 Resistor~
219 217 150 0 3 5
0 8 4 1
0
0 0 608 0
2 1k
-7 -14 7 -6
2 R1
-6 -14 8 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
972 0 0
2
44500.7 9
0
11
0 0 3 0 0 4096 0 0 0 10 0 2
341 144
368 144
2 0 4 0 0 4096 0 7 0 0 4 2
254 158
254 150
1 1 2 0 0 4224 0 2 7 0 0 4
254 199
254 202
254 202
254 194
1 2 4 0 0 4224 0 6 10 0 0 2
274 150
235 150
1 1 5 0 0 8320 0 3 8 0 0 3
178 67
178 75
200 75
1 3 6 0 0 4224 0 4 6 0 0 2
292 125
292 131
2 0 7 0 0 4096 0 8 0 0 11 2
236 75
254 75
1 1 8 0 0 8320 0 1 10 0 0 3
178 143
178 150
199 150
1 4 9 0 0 12416 0 5 6 0 0 4
292 167
292 168
292 168
292 157
2 5 3 0 0 8320 0 9 6 0 0 4
316 75
341 75
341 144
310 144
1 2 7 0 0 8320 0 9 6 0 0 4
280 75
254 75
254 138
274 138
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
283 177 308 201
287 181 303 197
2 -V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
283 91 308 115
287 95 303 111
2 +V
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
350 127 371 145
354 131 366 143
2 Vo
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
100 1 0.1 1e+06
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
4719804 1210432 100 100 0 0
0 0 0 0
11 334 172 404
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 5
1
339 75
0 3 0 0 1	0 10 0 0
4654234 8550464 100 100 0 0
77 66 377 156
400 74 800 322
377 66
77 66
377 66
377 156
0 0
0 0 0 0 0 0
12401 0
4 0.001 10
2
329 144
0 3 0 0 3	0 10 0 0
191 150
0 8 0 0 1	0 8 0 0
3540064 4356160 100 100 0 0
77 66 371 156
400 322 799 570
371 66
77 66
371 66
371 156
0 0
0 0 0 0 0 0
12403 0
4 0.3 5
1
334 144
0 2 0 0 3	0 10 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
