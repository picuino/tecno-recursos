CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 80 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
10
10 Op-Amp5:A~
219 291 144 0 5 11
0 4 3 6 7 5
0
0 0 64 0
6 OPAMP5
16 -25 58 -17
2 U1
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 26133460
88 0 0 0 1 1 0 0
1 U
7168 0 0
2
44500.7 0
0
2 +V
167 172 180 0 1 3
0 8
0
0 0 53856 0
2 5V
-8 -22 6 -14
3 Vi2
-9 -13 12 -5
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3171 0 0
2
5.89977e-315 0
0
2 +V
167 172 122 0 1 3
0 9
0
0 0 53856 0
2 5V
-8 -22 6 -14
3 Vi1
-9 -13 12 -5
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4139 0 0
2
5.89977e-315 5.26354e-315
0
2 +V
167 291 113 0 1 3
0 6
0
0 0 53344 0
3 15V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6435 0 0
2
5.89977e-315 5.32571e-315
0
2 +V
167 291 186 0 1 3
0 7
0
0 0 53344 180
4 -15V
-12 12 16 20
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5283 0 0
2
5.89977e-315 5.34643e-315
0
7 Ground~
168 255 254 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6874 0 0
2
5.89977e-315 5.3568e-315
0
9 Resistor~
219 255 228 0 3 5
0 2 3 -1
0
0 0 608 90
2 1k
8 0 22 8
2 RA
5 -4 19 4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 26134880
82 0 0 0 1 0 0 0
1 R
5305 0 0
2
44500.7 1
0
9 Resistor~
219 201 195 0 3 5
0 8 4 1
0
0 0 608 0
2 1k
-7 -14 7 -6
2 R2
-7 -13 7 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
34 0 0
2
5.89977e-315 5.36716e-315
0
9 Resistor~
219 298 204 0 2 5
0 3 5
0
0 0 608 0
2 2k
-7 -14 7 -6
2 RF
-7 6 7 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
969 0 0
2
5.89977e-315 5.38788e-315
0
9 Resistor~
219 201 138 0 3 5
0 9 4 1
0
0 0 608 0
2 1k
-7 -14 7 -6
2 R1
-7 -13 7 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8402 0 0
2
5.89977e-315 5.39306e-315
0
11
1 0 3 0 0 4112 0 9 0 0 6 2
280 204
255 204
1 0 4 0 0 4096 0 1 0 0 3 2
273 138
235 138
2 2 4 0 0 0 0 10 8 0 0 4
219 138
236 138
236 195
219 195
0 0 5 0 0 4096 0 0 0 5 0 2
337 144
366 144
2 5 5 0 0 8320 0 9 1 0 0 4
316 204
337 204
337 144
309 144
2 2 3 0 0 8320 0 1 7 0 0 3
273 150
255 150
255 210
1 1 2 0 0 4224 0 6 7 0 0 4
255 248
255 251
255 251
255 246
3 1 6 0 0 4224 0 1 4 0 0 2
291 131
291 122
1 4 7 0 0 4224 0 5 1 0 0 2
291 171
291 157
1 1 8 0 0 4224 0 2 8 0 0 3
172 189
172 195
183 195
1 1 9 0 0 4224 0 3 10 0 0 3
172 131
172 138
183 138
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
280 178 305 202
284 182 300 198
2 -V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
280 91 305 115
284 95 300 111
2 +V
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
349 125 370 143
353 129 365 141
2 Vo
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
100 1 0.1 1e+06
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2032918 1210432 100 100 0 0
0 0 0 0
486 365 647 435
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 10
1
334 144
0 2 0 0 3	0 12 0 0
2098462 8550464 100 100 0 0
77 66 377 156
400 74 800 322
377 66
77 66
377 66
377 156
0 0
0 0 0 0 0 0
12401 0
4 0.001 10
1
340 144
0 2 0 0 1	0 12 0 0
3540064 4356160 100 100 0 0
77 66 371 156
400 322 799 570
371 66
77 66
371 66
371 156
0 0
0 0 0 0 0 0
12403 0
4 0.3 5
1
334 144
0 2 0 0 3	0 12 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
