��  CCircuit��  CSerializeHack           ��  CPart�� 	 CGroupBox  D�T�             �  $ ��             �  D$ T�             �  $ $ �                           ���  CMotorEM�� 	 CTerminal  ��%        '�=� �>�C�Ƽ  �  ����     
  ��=� �>�C��<  �� 	 CMechTerm�j:IR��              P�    \              %     	 �j:IR��      P�    �$�        ��  D `  bK�6�>�j:IR��         ��433���j:IR��        ��  xy%      	          �          �  x�y�               �          �       �                    \             � �%     	        �            `$��         ��  D `  bK�6�>       �                       �        ��  �� ��          6��]���?(� !�C�?  �  ��)          X����>(� !�C��  �<�j;]����2u|�m�      �<    \             � �      	 <�j;]���      �<    ��         ��  D `  bK�6�><�j;]���+�t�a����[����<�j;]���+�t�a�����  x� y�                 �          �  xy)                           ��?( �                    \             �� ��      	 �?( �            `� �        ��  D `  bK�6�>�?( ��T�r��  f �)�?( ��T�r����  CBattery��  CDummyValue  �8�8    1.5V            �?      �? V �  �(�=         [�~���?��>���  �  ����     
  ��=� �  X�b�ɼ    �<��     $    ��   �   �"�  x8x8    1.5V            �?      �? V �  x(y=         ������@          �  x�y�        [�~���?��>��=    h<��     (    ��   �  �� 	 CPushMake��  CKey  �"�      +  �  �	        ������@          �  �       '�=� �            ��!�     .    ����    �� 
 CBattery9V"�  � H� H    9V            "@      �? V �  � 8� M                �          �  ` 8a M              "@            L L� �     3    ��   �  *�,�  � �� �      5  �  � ��              "@          �  � ��      	          �            � �� �     7    ����    �� 
 CVResistor��  CSlider  �i o�     "�  �� ��     100            Y@      �?    = �  �� ��        ���u "@�� !�C�?  �  t� ��         6��]���?�� !�C��    �� t�      >      ���   0�"�  �� ��     9V            "@      �? V �  �� ��            X����>(� !�C�?  �  x� y�         ���u "@�� !�C��    d� �h     B    ��   �  0�"�  � � � �     9V            "@      �? V �  � � � �                            �  X � Y �               "@            D � � h     F    ��   �  ��  CSPST��  CToggle  � @  d       I  �  � � � �              "@          �  � � � �                �            � b  �      L    ����P                  ���  CWire  ����      
 O�  ����     
 O�  �      O�  �� ��       O�  H�y�      O�  H8I�       O�  � 8I9      O�  � y     	 O�  �(�)      O�  �� �)       O�  �� ��       O�  H(y)       O�  H� I)        O�  � � I�        O�  � � y�       O�  x	      O�  xy)       O�  �(�)      O�  �(��       O�  x���      O�  ` a 9       O�  ` �       O�  X � � �       O�  x� y�        O�  x� ��       O�  X � Y �                      �                             R    P      W    T      Z    X      ^    [     $ a $ % % Q ( ` ( ) ) c . . _ / / R 3 V 3 4 d 4 7 7 e 8 8 W > h > ? ? Z B S B C g C F ] F G i G L L f M M ^  Q % P /  B Y U  V T 3 U 8  Y  S X ?  \  ] [ F \ M  ` . _ ( b $ a c ) b e 4 d 7 i L h C g > f G   D        �4s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 