CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
21 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
18
8 Op-Amp5~
219 405 100 0 5 11
0 7 3 6 5 3
0
0 0 64 0
5 UA741
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 1 0 0
1 U
317 0 0
2
5.90009e-315 5.30499e-315
0
2 +V
167 405 72 0 1 3
0 6
0
0 0 53344 0
3 15V
-11 -27 10 -19
2 V4
-7 -15 7 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3108 0 0
2
5.90009e-315 5.26354e-315
0
2 +V
167 405 133 0 1 3
0 5
0
0 0 53344 180
4 -15V
-13 12 15 20
2 V3
-5 0 9 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4299 0 0
2
5.90009e-315 0
0
7 Ground~
168 366 177 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9672 0 0
2
5.90009e-315 0
0
10 Capacitor~
219 343 106 0 2 5
0 4 7
0
0 0 576 0
6 0.02uF
-22 -18 20 -10
2 C4
-6 -20 8 -12
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7876 0 0
2
5.90009e-315 0
0
10 Capacitor~
219 304 106 0 2 5
0 8 4
0
0 0 576 0
6 0.02uF
-22 -18 20 -10
2 C3
-6 -20 8 -12
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6369 0 0
2
5.90009e-315 0
0
10 Capacitor~
219 190 26 0 2 5
0 9 8
0
0 0 576 0
6 0.02uF
-22 -18 20 -10
2 C2
-6 -20 8 -12
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9172 0 0
2
5.90009e-315 5.37752e-315
0
2 +V
167 253 139 0 1 3
0 11
0
0 0 53344 180
4 -15V
-13 12 15 20
2 V2
-5 0 9 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7100 0 0
2
5.90009e-315 5.36716e-315
0
2 +V
167 253 79 0 1 3
0 12
0
0 0 53344 0
3 15V
-11 -27 10 -19
2 V1
-7 -15 7 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3820 0 0
2
5.90009e-315 5.3568e-315
0
7 Ground~
168 114 176 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7678 0 0
2
5.90009e-315 5.34643e-315
0
7 Ground~
168 213 176 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
961 0 0
2
5.90009e-315 5.32571e-315
0
11 Signal Gen~
195 76 117 0 64 64
0 10 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 64 0
5 -1/1V
-18 -30 17 -22
2 Vi
-6 -33 8 -25
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 1 0 0
1 V
3178 0 0
2
5.90009e-315 5.30499e-315
0
10 Capacitor~
219 213 153 0 2 5
0 2 13
0
0 0 576 90
6 0.01uF
10 0 52 8
2 C1
13 -3 27 5
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3409 0 0
2
5.90009e-315 5.26354e-315
0
8 Op-Amp5~
219 253 106 0 5 11
0 13 8 12 11 8
0
0 0 64 0
5 UA741
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 1 0 0
1 U
3951 0 0
2
5.90009e-315 0
0
9 Resistor~
219 358 27 0 2 5
0 4 3
0
0 0 608 0
6 11.25k
-21 -14 21 -6
2 R4
-5 -13 9 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8885 0 0
2
5.90009e-315 0
0
9 Resistor~
219 366 145 0 3 5
0 2 7 -1
0
0 0 608 90
6 11.25k
-21 -14 21 -6
2 R3
4 -4 18 4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3780 0 0
2
5.90009e-315 0
0
9 Resistor~
219 135 112 0 2 5
0 10 9
0
0 0 608 0
6 11.25k
-21 -14 21 -6
2 R1
-4 -14 10 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9265 0 0
2
5.90009e-315 5.39306e-315
0
9 Resistor~
219 189 112 0 2 5
0 9 13
0
0 0 608 0
6 11.25k
-21 -14 21 -6
2 R2
-5 -13 9 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9442 0 0
2
5.90009e-315 5.38788e-315
0
21
1 1 0 0 0 0 0 12 17 0 0 2
107 112
117 112
2 0 3 0 0 4096 0 15 0 0 6 3
376 27
441 27
441 49
1 0 4 0 0 8320 0 15 0 0 10 3
340 27
323 27
323 106
1 4 5 0 0 4224 0 3 1 0 0 2
405 118
405 113
1 3 6 0 0 4224 0 2 1 0 0 2
405 81
405 87
2 5 3 0 0 12416 0 1 1 0 0 6
387 94
367 94
367 49
441 49
441 100
423 100
2 1 7 0 0 4224 0 0 1 9 0 4
366 106
395 106
395 106
387 106
1 1 2 0 0 4096 0 4 16 0 0 2
366 171
366 163
2 2 7 0 0 0 0 16 5 0 0 3
366 127
366 106
352 106
1 2 4 0 0 0 0 5 6 0 0 2
334 106
313 106
1 0 8 0 0 4096 0 6 0 0 18 3
295 106
282 106
282 105
1 1 2 0 0 0 0 11 13 0 0 2
213 170
213 162
2 0 8 0 0 4224 0 7 0 0 18 3
199 26
282 26
282 49
1 0 9 0 0 8320 0 7 0 0 15 3
181 26
166 26
166 112
2 1 9 0 0 0 0 17 18 0 0 2
153 112
171 112
1 4 11 0 0 4224 0 8 14 0 0 2
253 124
253 119
1 3 12 0 0 4224 0 9 14 0 0 2
253 88
253 93
2 5 8 0 0 0 0 14 14 0 0 6
235 100
212 100
212 49
282 49
282 106
271 106
1 2 2 0 0 4224 0 10 12 0 0 3
114 170
114 122
107 122
2 0 13 0 0 4224 0 13 0 0 21 2
213 144
213 112
2 1 13 0 0 0 0 18 14 0 0 4
207 112
236 112
236 112
235 112
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
61 76 88 100
66 80 82 96
2 Vi
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
413 75 450 99
423 83 439 99
2 Vo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
234 128 271 152
244 136 260 152
2 -V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
236 53 273 77
246 61 262 77
2 +V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
387 46 424 70
397 54 413 70
2 +V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
388 122 425 146
398 130 414 146
2 -V
0
9 0 0
0
0
2 V1
-0.7 -1.5 -0.02
0
0 0 0
100 0 10 10000
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2032608 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 5e-06 10
0
2163704 4421696 100 100 0 0
77 66 779 156
-4 333 798 572
545 66
779 66
779 73
779 151
0 0
0 0 0 0 0 0
12403 4
4 500 1000
1
369 149
0 3 0 0 3	0 22 0 0
6030466 4421696 100 100 0 0
77 66 767 156
-4 333 798 572
86 66
77 66
767 97
767 97
0 0
0 0 0 0 0 0
12401 0
4 20 0.5
1
324 112
0 5 0 0 3	0 22 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
