CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
21 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
10
8 Op-Amp5~
219 317 149 0 5 11
0 8 3 7 6 3
0
0 0 64 0
5 UA741
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 1 0 0
1 U
3472 0 0
2
44525.3 0
0
10 Capacitor~
219 277 198 0 2 5
0 2 8
0
0 0 576 90
6 0.01uF
10 0 52 8
2 C1
13 -3 27 5
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9998 0 0
2
44525.3 1
0
11 Signal Gen~
195 105 160 0 64 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162722
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 64 0
5 -1/1V
-18 -30 17 -22
2 Vi
-6 -33 8 -25
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 1 0 0
1 V
3536 0 0
2
44525.3 2
0
7 Ground~
168 277 225 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
44525.3 3
0
7 Ground~
168 136 225 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3835 0 0
2
44525.3 4
0
2 +V
167 317 122 0 1 3
0 7
0
0 0 53344 0
3 15V
-11 -27 10 -19
2 V1
-7 -15 7 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3670 0 0
2
44525.3 5
0
2 +V
167 317 182 0 1 3
0 6
0
0 0 53344 180
4 -15V
-13 12 15 20
2 V2
-5 0 9 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5616 0 0
2
44525.3 6
0
10 Capacitor~
219 245 70 0 2 5
0 4 3
0
0 0 576 0
6 0.02uF
-22 -18 20 -10
2 C2
-6 -20 8 -12
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9323 0 0
2
44525.3 7
0
9 Resistor~
219 239 155 0 2 5
0 4 8
0
0 0 608 0
6 11.25k
-21 -14 21 -6
2 R2
-5 -13 9 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
317 0 0
2
44525.3 8
0
9 Resistor~
219 173 155 0 2 5
0 5 4
0
0 0 608 0
6 11.25k
-21 -14 21 -6
2 R1
-4 -14 10 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3108 0 0
2
44525.3 9
0
11
1 1 2 0 0 4096 0 4 2 0 0 2
277 219
277 207
2 0 3 0 0 4224 0 8 0 0 8 3
254 70
375 70
375 92
1 0 4 0 0 8320 0 8 0 0 5 3
236 70
206 70
206 155
1 1 5 0 0 4224 0 10 3 0 0 2
155 155
136 155
2 1 4 0 0 0 0 10 9 0 0 2
191 155
221 155
1 4 6 0 0 4224 0 7 1 0 0 2
317 167
317 162
1 3 7 0 0 4224 0 6 1 0 0 2
317 131
317 136
2 5 3 0 0 0 0 1 1 0 0 6
299 143
276 143
276 92
375 92
375 149
335 149
1 2 2 0 0 4224 0 5 3 0 0 2
136 219
136 165
2 0 8 0 0 4096 0 2 0 0 11 2
277 189
277 155
2 1 8 0 0 4224 0 9 1 0 0 4
257 155
300 155
300 155
299 155
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
93 118 120 142
98 122 114 138
2 Vi
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
346 122 383 146
356 130 372 146
2 Vo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
298 171 335 195
308 179 324 195
2 -V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
300 96 337 120
310 104 326 120
2 +V
0
9 0 0
0
0
2 V1
-0.7 -1.5 -0.02
0
0 0 0
100 0 10 10000
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2032608 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 5e-06 10
0
2163704 4421696 100 100 0 0
77 66 779 156
-4 333 798 572
545 66
779 66
779 73
779 151
0 0
0 0 0 0 0 0
12403 4
4 500 1000
1
369 149
0 3 0 0 3	0 8 0 0
6030466 4421696 100 100 0 0
77 66 767 156
-4 333 798 572
86 66
77 66
767 97
767 97
0 0
0 0 0 0 0 0
12401 0
4 20 0.5
1
324 112
0 5 0 0 3	0 12 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
