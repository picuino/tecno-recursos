CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
5
2 +V
167 166 75 0 1 3
0 2
0
0 0 53856 0
3 10V
-11 -22 10 -14
3 Vi2
-10 -15 11 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
5.89601e-315 0
0
2 +V
167 134 93 0 1 3
0 4
0
0 0 53856 0
3 10V
-11 -22 10 -14
3 Vi1
-10 -15 11 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
44269.4 0
0
2 +V
167 243 76 0 1 3
0 5
0
0 0 53344 0
3 15V
-10 -14 11 -6
3 Vi4
-10 -24 11 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3536 0 0
2
44269.4 1
0
2 +V
167 243 160 0 1 3
0 6
0
0 0 53344 180
4 -15V
-14 -1 14 7
3 Vi3
-10 0 11 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4597 0 0
2
44269.4 2
0
8 Op-Amp5~
219 243 114 0 5 11
0 4 2 5 6 3
0
0 0 64 0
5 LF353
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 589828
88 0 0 0 2 1 1 0
1 U
3835 0 0
2
44269.4 3
0
5
1 2 2 0 0 8320 0 1 5 0 0 3
166 84
166 108
225 108
5 0 3 0 0 4224 0 5 0 0 0 2
261 114
305 114
1 1 4 0 0 8320 0 2 5 0 0 3
134 102
134 120
225 120
3 1 5 0 0 4224 0 5 3 0 0 2
243 101
243 85
1 4 6 0 0 4224 0 4 5 0 0 2
243 145
243 127
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
231 156 256 180
235 160 251 176
2 -V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
231 50 256 74
235 54 251 70
2 +V
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
287 96 308 114
291 100 303 112
2 Vo
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.0175 7e-05 7e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2425688 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 10
0
2491180 8550464 100 100 0 0
77 66 767 156
0 322 800 570
472 66
77 66
767 66
767 156
0 0
0 0 0 0 0 0
12401 0
4 0.01 10
2
116 108
0 7 0 0 1	0 6 0 0
272 114
0 3 0 0 1	0 6 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
