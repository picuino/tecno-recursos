��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  AR    S6      �  � �     S5      �  A R     S4      �  A�R�    S3      �  � �� �    S2      �  A �R �    S1      �  � 9� G    S1      �  A�R�    S6      �  � �� �    S5      �  A �R �    S4      �  AiRw    S3      �  � i� w    S2      �  A iR w    S1      �  Y� j�     S6      �  � � � �     S5      �  YY jg     S4      �  � i � w     S3      �  Q y b �     S2        � � � �     ���  CSPDT��  CToggle  8�X          �� 	 CTerminal  (�=�                          �  T�i�     #                     �  T�i�               �            <�T�            ��    ��  8xX�      #   �  (h=i     "                     �  Tpiq               �          �  T`ia     !          �            <\Tt     %      ��    ��  � ��        (   �  � �� �                           �  � �� �     "                     �  � �� �     #                       � �� �     *      ��    ��  � x� �      -   �  � h� i                           �  � p� q     !          �          �  � `� a                            � \� t     /      ��    ��  CBulb�  $@9A                          �  � @A                             4$L    4    ��      ��  CBattery��  CValue  t '� 5    9V         "@      �? V �  h @} A             "@          �  � @� A                            | 4� L    :    ��      ��  8 �X        <   �  ( �= �               �          �  T �i �             "@          �  T �i �                            < �T �     >      ��    ��  8 xX �      A   �  ( h= i             "@          �  T pi q               �          �  T `i a             "@            < \T t     C      ��    ��  8�X�      F   �  (�=�                          �  T�i�               �          �  T�i�                            <�T�     H      ��    ��  8HXh      K   �  (8=9                          �  T@iA                          �  T0i1                            <,TD     M      ��    ��  � �� �      P   �  � �� �               �          �  � �� �               �          �  � �� �                            � �� �     R      ��    ��  � H� h      U   �  � 8� 9                          �  � @� A               �          �  � 0� 1                            � ,� D     W      ��    2��  $9               �          �  �                             $    [    ��      6�8�  t ��     9V         "@      �? V �  h }              "@          �  � �                            | �     _    ��      ��  8 �X �      a   �  ( �= �             "@          �  T �i �               �          �  T �i �             "@            < �T �     c      ��    ��  8 HX h      f   �  ( 8= 9             "@          �  T @i A             "@          �  T 0i 1             "@            < ,T D     h      ��    ��  CDPDT�  H X h x       l   �  8 ( M )                �          �  8 H M I                           �  d P y Q                �          �  d @ y A                           �  d 0 y 1                           �  d   y !                             L  d T      n      �� ,   ��  CSPST�  � � �       u   �  � � � �                �          �  � � � �              "@            � � � �      w      ��    6�8�  � <�     9V         "@      �? V �  � �              "@          �  4� I�      
         �            � 4�     {    ��      2��  �� ��                 �          �  �� ��      
          �            �� ��      ~    ��      ��  � �  �       �   �  � � � �                           �  � � �      	                     �  � � �                �            � | � �      �      ��    ��  P� p�       �   �  l� ��                �          �  @� U�                           �  @� U�      	                       T| l�     �      ��    ��  P8 pX       �   �  l( �)                           �  @  U!                           �  @0 U1                             T l4     �      ��    ��  � H  h       �   �  � 8 � 9                �          �  � @ A                �          �  � 0 1                             � , � D      �      ��      � � � �     ���  CWire�� 
 CCrossOver  � ��        � ��     # ����  � ��         h�      " ��  ��      # ����  f�l�        �y�     # ����  f�l�      ��  f�l�        hpi�       ����  v�|�        x�y�      # ����  v�|�      ��  f�l�        (���      ��  h�y�     # ��  hPia      ! ��  � PiQ     ! ����  � \� d        � P� q      ! ����  � \� d        � `� a      ��  � p� q     ! ��  h `� a      ����  ~ �� �        � `� �       ��  h �� �      ����  ~ �� �      ��  � �� �        h �� �      ��  h pi �       ��  ( �i �      ��  ( �) �       ��  h �i �       ����  � �� �        � h� �        ��  � `� �       ��  � h� i       ��  � �� �       ��  � ��     " ��   h)i     " ��  8@�A      ��  ���A       ��  (�)�       ��   h) i      ��   h A       ��   @i A      ��  � @� A       ��  h @i y       ��  ( xi y      ��  ( x) �       ��  h �y �      ��  x 0y �       ��  h 0y 1      ��  h �� �      ��  � �� �       ��  � �� �      ��  � x� �       ��  � x� y      ��  � 8� y       ��  � 0)1      ��  (0)9       ��  � @� A      ��  � @� �       ��  � �� �      ��  (x)�       ��  (xiy      ��  h@iy       ��  h0y1      ��  x0y�       ��  h�y�      ��   i       ��   8        ��   8) 9      ��  h�y�      ��  x�y       ��  8y      ��  � �       ��  �( �)       ��  �( �q        ��  @p �q       ��  @p A�        ��   � � �       ��   (  �        ��   ( 9 )       ��  � 8 � 9       ��  � 8 � Q        ����  � L � T       ��  � L � T         x P � Q       ����  � L � T         �   � �        ����  � L � T         � 0 � �        ��  x   � !       ��  x @ � A       ����  � , � 4         �   � A        ����  � , � 4         x 0 � 1       ��  ( � � �       ��  ( H 9 I       ��  ( H ) �        ��  � � 	�       ��  H� ��      
 ��  �� ��        ��  �� ��       ��  @ A       ��  @ �        ��  � �       ��  �   A!       ��  � � � �       ��  � A�      	 ��  0 A1         � � � �     �  � � � �       � � � �       �   ! ! � " " � % � % & & � ' ' � * � * + + � , , � / � / 0 0 � 1 1 � 4 4 � 5 � 5 : � : ; ; � > � > ? ? � @ @ � C � C D D � E E � H � H I I � J J � M � M N N � O O � R � R S S � T T � W � W X X � Y Y � [ [ � \ � \ _ � _ ` ` � c � c d d � e e � h � h i i � j j � n � n o � o p p � q q � r r � s s � w � w x x � { � { | | � ~  ~   � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � , � � � � � � � � � � � � � � � & " � � � � � � � � � � ! � � ' � � � � � � � � 1 � 0 � E � � � � � ? � � � � � � � D � � � � > � @ � � � � � � � / � * + � � % 4 � � � �   � C � � � : ; 5 i � � � � c e � � � j � d � � � � R � T � � W � Y � � M X � � � S � � H � � N � O � � � J � � _ � � � h I � � � [ � ` \ � � � � � � � � � w � � � n � � � � � � � � p � � � � � � � s � q � � � � � � � r � � � � o � � x { |  ~ �  � � � � � � � � � �  $ 7         �$s�        @     +        @            @    "V  (      X�                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 