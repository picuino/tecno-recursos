��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  	    S2      �  	� �     S1      �  ����    L2      �  �Y�g    L1      �  Y� i�     L1      �  � Q � _     S1      �  � � � �     S2                    ���  CBattery��  CValue  � �     9V         "@      �? V �� 	 CTerminal  �( )              "@          �  �( �)                             � �4         ��      �� 	 CRailThru�   ( 5)       e       "@          �  $( 9)              "@            "$ 6,          ����    ��   H 5I        d                   �  $H 9I                             "D 6L          ����    ��   � 5�       d        �          �  $� 9�                             "� 6�          ����    ��  CSPDT��  CToggle  ��(      "   �  �� 	�                �          �  �� ��                �          �  � �                            �� �    %      ��    ��   (5)      d                   �  $(9)                            "$6,     )    ����    ��    5      d        �          �  $ 9                            "� 6     ,    ����    ��   � 5�       d        �          �  $� 9�                             "� 6�      /    ����    ��   � 5�       d                   �  $� 9�                             "� 6�      2    ����    !�#�  �� ��       4   �  �� 	�                �          �  �� ��                �          �  �� ��                             �| ��     6      ��    ��   h 5i       d        �          �  $h 9i                             "d 6l      :    ����    ��   H5I     
 d        �          �  $H9I                            "D6L     =    ����    ��  CBulb�  �HI     
          �          �  �H�I               �            �<�T    A    ��      ��   h5i      d        �          �  $h9i     	                       "d6l     D    ����    ��   �5�      d        �          �  $�9�                            "�6�     G    ����    ?��  ���               �          �  ����               �            �|��    J    ��      ��   �5�      d        �          �  $�9�                            "�6�     M    ����    ��   � 3 �     9V(          "@      �? V �  @ � A �               "@          �  @ � A �                             4 � L �      Q    ��      ?��  H� I�                 �          �  H� I�                             <� T�      T    ��      ��  CSPST#�  � 0 � P       W   �  � ( � )              "@          �  � ( � )                �            � $ � ,      Y      ��    V�#�  � � � �       [   �  � � � �              "@          �  � � � �                �            � | � �      ]      ��                  ���  CWire   ( !)       `�  �H !I        `�  �( �I         `�  �( �)        `�  �� ��       `�  �� ��        `�  �� !�       `�  � �       `�  �        `�   !      `�  �(!)      `�  � �)       `�  � �      `�  �� ��       `�  �� ��        `�  �� !�       `�  � !�       `�  � �        `�  � �       `�  �h !i       `�  �h ��        `�  �� ��       `�  H!I     
 `�  �h!i      `�  �H�i       `�  �H�I      `�  ����      `�  ����       `�  ��!�      `�  �!�      `�  @ � A �        `�  @ � I�       `�  H� I�        `�  @ ( A �        `�  � � � �       `�  � ( � �        `�  � ( � )       `�  � � � �       `�  � ( � �        `�  @ ( � )       `�  � ( � )       `�  � ( I)       `�  H( I�                      �                              a  d  a      b      g        % % h & e & ' m ' k ) * *   j , - -   q / 0 0   p 2 3 3   6 6 s 7 v 7 8 n 8 t : ; ;   w = > >   A A w B z B x D E E   } G H H   J J ~ K { K ~ M N N   Q � Q R R  T � T U U � Y � Y Z Z � ] � ] ^ ^ �   c  d b c  f & g e f  % i h j i , l ) m k l ' o 8 n p o 2 r / s q 6 r u : t v u 7 A = y D z x y B | K { } | G J M R �  � U � � Q ^ � � � Z � � ] � � � � � Y � � � T            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 