CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
21 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
12
2 +V
167 318 194 0 1 3
0 6
0
0 0 53344 180
4 -15V
-13 12 15 20
2 V2
-5 0 9 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3674 0 0
2
44525.5 2
0
2 +V
167 318 134 0 1 3
0 7
0
0 0 53344 0
3 15V
-11 -27 10 -19
2 V1
-7 -15 7 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5697 0 0
2
44525.5 1
0
8 Op-Amp5~
219 318 161 0 5 11
0 8 3 7 6 3
0
0 0 64 0
5 UA741
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 1 0 0
1 U
3805 0 0
2
44525.5 0
0
7 Ground~
168 206 216 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5219 0 0
2
44525.5 0
0
9 Resistor~
219 206 187 0 1 5
0 0
0
0 0 608 90
2 1k
8 0 22 8
2 Rr
4 -7 18 1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 39066004
82 0 0 0 1 0 0 0
1 R
3795 0 0
2
44525.5 0
0
10 Capacitor~
219 242 155 0 2 5
0 2 8
0
0 0 576 180
6 0.01uF
10 0 52 8
2 C1
-7 -18 7 -10
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3637 0 0
2
5.90009e-315 5.26354e-315
0
11 Signal Gen~
195 113 160 0 64 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162722
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 64 0
5 -1/1V
-18 -30 17 -22
2 Vi
-6 -33 8 -25
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 1 0 0
1 V
3226 0 0
2
5.90009e-315 5.30499e-315
0
7 Ground~
168 277 216 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6966 0 0
2
5.90009e-315 5.32571e-315
0
7 Ground~
168 150 215 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9796 0 0
2
5.90009e-315 5.34643e-315
0
10 Capacitor~
219 245 70 0 2 5
0 4 3
0
0 0 576 0
6 0.02uF
-22 -18 20 -10
2 C2
-6 -20 8 -12
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5952 0 0
2
5.90009e-315 5.37752e-315
0
9 Resistor~
219 316 99 0 2 5
0 4 8
0
0 0 608 0
6 11.25k
-21 -14 21 -6
2 R2
-5 -13 9 -5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3649 0 0
2
5.90009e-315 5.38788e-315
0
9 Resistor~
219 173 155 0 2 5
0 5 4
0
0 0 608 0
6 11.25k
-21 -14 21 -6
2 R1
-4 -14 10 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3716 0 0
2
5.90009e-315 5.39306e-315
0
13
1 1 0 0 0 0 0 3 8 0 0 3
300 167
277 167
277 210
2 0 0 0 0 0 0 11 0 0 10 2
334 99
369 99
1 0 0 0 0 0 0 11 0 0 4 3
298 99
277 99
277 155
2 1 0 0 0 0 0 3 6 0 0 2
300 155
251 155
1 4 6 0 0 0 0 1 3 0 0 2
318 179
318 174
1 3 7 0 0 0 0 2 3 0 0 2
318 143
318 148
2 0 0 0 0 0 0 6 0 0 9 2
233 155
206 155
1 1 0 0 0 0 0 4 5 0 0 4
206 210
206 212
206 212
206 205
2 0 0 0 0 0 0 5 0 0 11 2
206 169
206 155
2 5 3 0 0 4224 0 10 3 0 0 4
254 70
369 70
369 161
336 161
1 2 4 0 0 8320 0 10 12 0 0 4
236 70
206 70
206 155
191 155
1 1 5 0 0 4224 0 12 7 0 0 2
155 155
144 155
1 2 2 0 0 4240 0 9 7 0 0 3
150 209
150 165
144 165
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
299 183 336 207
309 191 325 207
2 -V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
301 108 338 132
311 116 327 132
2 +V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
339 137 376 161
349 145 365 161
2 Vo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
101 118 128 142
106 122 122 138
2 Vi
0
9 0 0
0
0
2 V1
-0.7 -1.5 -0.02
0
0 0 0
100 0 10 10000
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2032608 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 5e-06 10
0
2163704 4421696 100 100 0 0
77 66 779 156
-4 333 798 572
545 66
779 66
779 73
779 151
0 0
0 0 0 0 0 0
12403 4
4 500 1000
1
369 149
0 3 0 0 3	0 14 0 0
6030466 4421696 100 100 0 0
77 66 767 156
-4 333 798 572
86 66
77 66
767 97
767 97
0 0
0 0 0 0 0 0
12401 0
4 20 0.5
1
324 112
0 5 0 0 3	0 14 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
