��  CCircuit��  CSerializeHack           ��  CPart  0   0       ��� 
 CPushBreak��  CKey  � � .      	   �� 	 CTerminal  p � 	             "@
ףp=
�?  �  � � 	             "@
ףp=
��    � �            ��    ��  CBattery��  CValue   1; ?    9V(          "@      �? V �  H I -              "@
ףp=
��  �  H DI Y               
ףp=
�?    < ,T D         ��      ��  CBulb�  � � -              "@
ףp=
�?  �  � D� Y                
ףp=
��    � ,� D       
 ��      �� 	 CPushMake
�  � � � �          �  p � � �              "@          �  � � � �                �            � � � �            ��    ��   A ; O     9V(          "@      �? V �  H ( I =               "@          �  H T I i                             < < T T           ��      ��  � ( � =                 �          �  � T � i                              � < � T      #    ��      ��  CSPST��  CToggle  �   � @       &   �  p  �               "@          �  �  �                 �            �  �       )      ��    ��  � � � �                 �          �  � � � �                �            � � � �      ,    ��      ��   � ; �     9V(          "@      �? V �  H � I �               "@          �  H � I �               �            < � T �      0    ��        0   0       ���  CWire  H I        3�  H q 	      3�  � �        3�  � � 	      3�  H X� Y      3�  H � I �        3�  H � q �       3�  � � � �        3�  � � � �       3�  H  q        3�  H  I )        3�  H h � i        3�  �  � )        3�  �  �        3�  H � � �         0   0       �  0   0         0   0        5    7  4    8  6    8  :    <   >   ! ! ? # @ # $ $ ? ) = ) * * A , ; , - - B 0 9 0 1 1 B 5  4  7   6   : 0 9  < ,  ; > ) =   ! $ A # * @ 1 -  	          �5s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 