��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  Aq Q     L2      �  � q �      L1      �  	9 G     S2      �  � 9 � G     S1      �  �Y	g    L1      �  ��	�    L2      �  � *�     S1      �  *    S2                    ���  CBulb�� 	 CTerminal  0X 1m                 �          �  0� 1�                �            $l <�          ��      ��  � X � m                 �          �  � � � �                �            � l � �          ��      ��  CSPST��  CToggle  � 0  P          �  � ( � )                �          �  � ( )                �            � $ � ,            ��    ��  h 0 � P          �  X ( m )              "@          �  � ( � )                �            l $ � ,      !      ��    �� 	 CRailThru�  0�E�      d                   �  4�I�               �            2�F�     %    ����    ��  �!�                          �  ����               �            �|�    (    ��      #��  0�E�      d        �          �  4�I�                            2�F�     +    ����    #��  0hEi      d        �          �  4hIi                            2dFl     .    ����    ��  H!I               �          �  �H�I               �            �<T    1    ��      #��  0HEI      d        �          �  4HII                            2DFL     4    ����    #��  0h Ei       d        �          �  4h Ii                             2d Fl      7    ����    ��  CSPDT�  �� �       :   �  � �                �          �  �� ��                �          �  �� ��                             �| �     <      ��    #��  0� E�       d                   �  4� I�                             2� F�      @    ����    #��  0� E�       d        �          �  4� I�                             2� F�      C    ����    #��  0 E      d        �          �  4 I                            2� F     F    ����    #��  0(E)      d                   �  4(I)                            2$F,     I    ����    9��  �(      K   �  � �                �          �  �� ��      	          �          �  � �                            ��     M      ��    #��  0� E�      	 d        �          �  4� I�      
                       2� F�      Q    ����    #��  0H EI        d                   �  4H II                             2D FL      T    ����    #��  0( E)       e       "@          �  4( I)              "@            2$ F,      W    ����    ��  CBattery��  CValue  �      9V         "@      �? V �  �( )              "@          �  �( �)                             � �4     ]    ��      Y�[�   Q 3 _     9V(          "@      �? V �  @ 8 A M               "@          �  @ d A y                �            4 L L d      a    ��                    ���  CWire  0( 1Y        d�  ( 1)       d�  � ( � Y        d�  � ( � )       d�  � ( � )       d�  @ x A �        d�  @ � � �       d�  � � 1�       d�  @ ( A 9        d�  @ ( Y )       d�   �1�      d�  ��1�      d�  ����       d�  ����      d�  �H�I      d�  �H�i       d�  �h1i      d�   H1I      d�  �� ��       d�  �h ��        d�  �h 1i       d�  � )�       d�  (� )�        d�  (� 1�       d�  �� 1�       d�  �� ��        d�  �� ��       d�  � �      d�  � �)       d�  �(1)      d�  ( 1      d�  (� )       d�  � )�       d�  �� 1�      	 d�  �� ��       	 d�  �� ��      	 d�  �( �)        d�  �( �I         d�  �H 1I        d�  ( 1)                     �                             e    l  g    l  i    f ! n ! " " h o % & &   ( ( o ) r ) p + , ,   u . / /   1 1 v 2 s 2 v 4 5 5   y 7 8 8   < < z = w = >  > } @ A A   | C D D   � F G G   � I J J   M M � N � N O � O � Q R R   � T U U   � W X X   ] ] � ^ � ^ a m a b b j f   e i  " g h  b k j  k  n a m ! ( % q + r p q ) t 2 s u t . 1 4 x = y w x 7 < { z | { C ~ @  } ~ > � O � � � I � F � � M � � Q � � � N � ^ � � � T ] W   Z         �%s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 