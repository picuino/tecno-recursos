��  CCircuit��  CSerializeHack           ��  CPart  � � � �     ���  CDPDT��  CToggle  H P h p       	   �� 	 CTerminal  8   M !                           �  8 @ M A                           �  d H y I                �          �  d 8 y 9      	          �          �  d ( y )                           �  d  y       	          �            L  d L            �� ,   ��  CSPST
�  � � �           �  � � � �                           �  � � � �      
        "@            � � � �            ��    ��  CBattery��  CValue  � <�     9V         "@      �? V �  � �      
        "@          �  4� I�                             � 4�         ��      ��  CBulb�  �� ��                 �          �  �� ��                              �� ��           ��      ��  CSPDT
�  � �  �       #   �  � � � �                           �  � � �                           �  � x y                �            � t � �      %      ��    "�
�  P� p�       (   �  l� ��                �          �  @x Uy                           �  @� U�                             Tt l�     *      ��    "�
�  P0 pP       -   �  l  �!                           �  @ U                           �  @( U)                             T l,     /      ��    "�
�  � @  `       2   �  � 0 � 1                �          �  � 8 9                �          �  � ( )                             � $ � <      4      ��      � � � �     ���  CWire   � � �       8�      �        8�     9 !       8�  � 0 � 1       8�  � 0 � I        8��� 
 CCrossOver  � D � L       ?�  � D � L         x H � I       8�?�  � D � L         �  � �        8�?�  � D � L         � ( � �        8�  x  �       	 8�  x 8 � 9      	 8�?�  � $ � ,         �  � 9       	 8�?�  � $ � ,         x ( � )       8�  ( � � �       8�  ( @ 9 A       8�  ( @ ) �        8�  � � 	�      
 8�  H� ��        8�  �� ��        8�  �� ��       8�  8 9       8�  8 y        8�  x y       8�  @X Ay        8�  @X �Y       8�  �  �Y        8�  �  A       8�  � � � �       8�  � A�       8�  ( A)         � � � �     �  � � � �       � � � �      ;   M    >   G   J   F  9    O  O    P   Q   ! ! P % Z % & & [ ' ' U * * R + V + , [ , / / X 0 Y 0 1 \ 1 4 < 4 5 5 S 6 6 \ :  ; 9 :  = 4 < > > C > E  = B @ Y Z D A J L  H  H H K F G J I  D N D N  M L    ! R   * Q 5 T S U ' T W + V X / W B 0 B % & , 6 1            �%s�        @     +        @            @    "V  (      X�                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 