CircuitMaker Text
5.6
Probes: 2
U1B_7
Transient Analysis
0 593 193 65280
U1B_7
AC Analysis
0 597 193 8421376
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 361
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
46 C:\Archivos de programa\CircuitMaker 6\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1446 465
144179218 0
0
6 Title:
5 Name:
0
0
0
19
10 Polar Cap~
219 324 36 0 2 5
0 10 11
0
0 0 592 180
5 0.1uF
-22 -18 13 -10
2 C2
-10 -20 4 -12
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9281 0 0
2
44525.6 0
0
10 Polar Cap~
219 254 179 0 2 5
0 12 11
0
0 0 592 180
5 0.1uF
-22 -18 13 -10
2 C1
-11 -20 3 -12
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8464 0 0
2
44525.6 1
0
7 Ground~
168 508 261 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7168 0 0
2
5.89939e-315 0
0
2 +V
167 535 260 0 1 3
0 4
0
0 0 53872 180
4 -10V
3 -2 31 6
2 V4
-6 1 8 9
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3171 0 0
2
5.89939e-315 5.26354e-315
0
2 +V
167 536 137 0 1 3
0 5
0
0 0 53872 0
3 10V
-11 -22 10 -14
2 V3
-5 -17 9 -9
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4139 0 0
2
5.89939e-315 5.30499e-315
0
2 +V
167 325 249 0 1 3
0 6
0
0 0 53872 180
4 -10V
3 -2 31 6
2 V2
-7 2 7 10
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6435 0 0
2
5.89939e-315 5.32571e-315
0
2 +V
167 325 138 0 1 3
0 7
0
0 0 53872 0
3 10V
-11 -22 10 -14
2 V1
-7 -17 7 -9
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5283 0 0
2
5.89939e-315 5.34643e-315
0
7 Ground~
168 93 233 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6874 0 0
2
5.89939e-315 5.3568e-315
0
11 Signal Gen~
195 46 184 0 19 64
0 9 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 Vi
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5305 0 0
2
5.89939e-315 5.36716e-315
0
7 Ground~
168 285 239 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
34 0 0
2
5.89939e-315 5.37752e-315
0
7 Ground~
168 212 277 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
969 0 0
2
5.89939e-315 5.38788e-315
0
8 Op-Amp5~
219 535 192 0 5 11
0 2 3 5 4 8
0
0 0 80 0
5 LF353
15 -25 50 -17
3 U1B
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 0 2 2 1 0
1 U
8402 0 0
2
5.89939e-315 5.39306e-315
0
8 Op-Amp5~
219 324 186 0 5 11
0 2 12 7 6 10
0
0 0 80 0
5 LF353
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 589827
88 0 0 0 2 1 1 0
1 U
3751 0 0
2
5.89939e-315 5.39824e-315
0
9 Resistor~
219 537 90 0 2 5
0 3 8
0
0 0 624 0
3 10k
-10 -14 11 -6
2 R5
-6 -16 8 -8
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4292 0 0
2
5.89939e-315 5.40342e-315
0
9 Resistor~
219 451 235 0 2 5
0 9 3
0
0 0 624 0
3 10k
-10 -14 11 -6
2 R4
-7 -15 7 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6118 0 0
2
5.89939e-315 5.4086e-315
0
9 Resistor~
219 450 186 0 2 5
0 10 3
0
0 0 624 0
3 10k
-10 -14 11 -6
2 R3
-7 -17 7 -9
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
34 0 0
2
5.89939e-315 5.41378e-315
0
9 Resistor~
219 212 237 0 3 5
0 2 11 -1
0
0 0 624 90
4 1332
6 1 34 9
2 Rr
-21 -2 -7 6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6357 0 0
2
5.89939e-315 5.41896e-315
0
9 Resistor~
219 160 179 0 2 5
0 9 11
0
0 0 624 0
6 265166
-21 -14 21 -6
2 R1
-6 -15 8 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
319 0 0
2
5.89939e-315 5.42414e-315
0
9 Resistor~
219 322 87 0 2 5
0 12 10
0
0 0 624 0
6 530333
-21 -14 21 -6
2 R2
-6 -14 8 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3976 0 0
2
5.89939e-315 5.42933e-315
0
22
1 1 2 0 0 4224 0 3 12 0 0 4
508 255
508 197
517 197
517 198
2 0 3 0 0 8192 0 15 0 0 8 3
469 235
486 235
486 185
1 4 4 0 0 4224 0 4 12 0 0 2
535 245
535 205
1 3 5 0 0 4224 0 5 12 0 0 3
536 146
536 179
535 179
1 4 6 0 0 4224 0 6 13 0 0 3
325 234
325 199
324 199
1 3 7 0 0 4224 0 7 13 0 0 3
325 147
325 173
324 173
2 5 8 0 0 8320 0 14 12 0 0 4
555 90
620 90
620 192
553 192
0 1 3 0 0 4224 0 0 14 10 0 3
486 186
486 90
519 90
0 1 9 0 0 8320 0 0 15 13 0 5
112 179
112 351
398 351
398 235
433 235
2 2 3 0 0 0 0 16 12 0 0 2
468 186
517 186
1 0 10 0 0 4096 0 16 0 0 21 2
432 186
400 186
1 2 2 0 0 0 0 8 9 0 0 3
93 227
93 189
77 189
1 1 9 0 0 0 0 9 18 0 0 2
77 179
142 179
1 1 2 0 0 0 0 10 13 0 0 3
285 233
285 192
306 192
1 1 2 0 0 0 0 11 17 0 0 2
212 271
212 255
2 0 11 0 0 4096 0 17 0 0 17 2
212 219
212 179
2 0 11 0 0 0 0 18 0 0 19 4
178 179
212 179
212 178
213 178
1 0 12 0 0 4096 0 2 0 0 22 3
261 179
286 179
286 180
2 2 11 0 0 8320 0 1 2 0 0 4
314 36
213 36
213 179
244 179
0 1 10 0 0 8192 0 0 1 21 0 3
400 87
400 36
331 36
2 5 10 0 0 8320 0 19 13 0 0 4
340 87
400 87
400 186
342 186
2 1 12 0 0 8320 0 13 19 0 0 4
306 180
286 180
286 87
304 87
0
0
2073 0 1
0
0
0
0 0 0
0
0 0 0
10000 0 1 1000
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
4654008 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 5
0
4391674 8550464 100 100 0 0
77 66 647 246
680 74 1360 406
647 66
77 66
647 66
647 246
0 0
0 0 0 0 0 0
12401 0
4 0.001 5
1
112 179
0 9 0 0 1	0 9 0 0
1311754 4356160 100 100 0 0
77 66 647 246
680 406 1360 738
647 66
77 66
647 67
647 246
0 0
0 0 0 0 0 0
12401 0
4 30 50
1
382 186
0 11 0 0 3	0 21 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
