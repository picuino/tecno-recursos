CircuitMaker Text
5.6
Probes: 1
RL_2
Transient Analysis
0 305 74 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1446 465
9961490 0
0
6 Title:
5 Name:
0
0
0
6
10 FW Bridge~
219 254 115 0 4 9
0 2 5 3 4
0
0 0 80 0
6 BRIDGE
-17 -50 25 -42
2 D2
-4 -60 10 -52
0
0
17 %D %1 %2 %3 %4 %S
0
0
0
9

0 1 2 3 4 1 2 3 4 0
88 0 0 256 0 0 0 0
1 D
9424 0 0
2
44470.7 0
0
7 Ground~
168 318 153 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9968 0 0
2
5.90002e-315 0
0
7 Ground~
168 142 152 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9281 0 0
2
5.90002e-315 0
0
7 Trans1~
219 171 110 0 4 9
0 6 2 5 4
0
0 0 592 0
5 10TO1
-17 -31 18 -23
2 T1
-6 -49 8 -41
0
0
17 %D %1 %2 %3 %4 %S
0
24 alias:XTRANS {RATIO=0.1}
0
9

0 1 2 3 4 1 2 3 4 0
88 0 0 0 1 0 0 0
1 T
8464 0 0
2
5.90002e-315 0
0
11 Signal Gen~
195 87 110 0 19 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1114636288 0 1120403456
20
1 60 0 100 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 592 0
9 -100/100V
-32 -30 31 -22
2 V1
-8 -31 6 -23
0
0
38 %D %1 %2 DC 0 SIN(0 100 60 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7168 0 0
2
5.90002e-315 0
0
9 Resistor~
219 318 116 0 3 5
0 2 3 -1
0
0 0 624 90
2 1k
8 0 22 8
2 RL
-18 -4 -4 4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 103767272
82 0 0 0 1 0 0 0
1 R
3171 0 0
2
5.90002e-315 0
0
8
1 0 2 0 0 4096 0 6 0 0 2 2
318 134
318 141
1 1 2 0 0 12416 0 1 2 0 0 7
224 111
216 111
216 161
295 161
295 141
318 141
318 147
3 2 3 0 0 8320 0 1 6 0 0 5
288 111
295 111
295 72
318 72
318 98
4 4 4 0 0 12416 0 4 1 0 0 5
189 127
198 127
198 149
256 149
256 143
3 2 5 0 0 12416 0 4 1 0 0 5
189 93
198 93
198 72
256 72
256 79
1 0 2 0 0 0 0 3 0 0 7 2
142 146
142 127
2 2 2 0 0 0 0 5 4 0 0 4
118 115
125 115
125 127
153 127
1 1 6 0 0 12416 0 5 4 0 0 4
118 105
125 105
125 93
153 93
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
320 105 347 129
325 109 341 125
2 Vo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
145 67 172 91
150 71 166 87
2 N1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
172 67 199 91
177 71 193 87
2 N2
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.0833333 0.000333333 0.000333333
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1705266 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 10
1
335 144
0 2 0 0 3	0 9 0 0
1967280 8550464 100 100 0 0
77 66 767 156
0 322 800 570
767 66
77 66
767 66
767 156
0 0
0 0 0 0 0 0
12385 0
4 1e-06 10
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
