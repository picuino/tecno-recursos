CircuitMaker Text
5.6
Probes: 2
V3_1
Transient Analysis
0 201 137 4227327
U1A_1
Transient Analysis
1 356 145 8421376
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 361
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1446 465
9961490 0
0
6 Title:
5 Name:
0
0
0
8
7 Ground~
168 206 165 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3440 0 0
2
5.90006e-315 0
0
11 Signal Gen~
195 158 143 0 19 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
5 -1/1V
-18 -30 17 -22
2 V3
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6263 0 0
2
5.90006e-315 5.26354e-315
0
2 +V
167 292 184 0 1 3
0 6
0
0 0 53600 180
4 -15V
7 -10 35 -2
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4900 0 0
2
5.90006e-315 5.30499e-315
0
2 +V
167 292 109 0 1 3
0 7
0
0 0 53600 0
3 15V
5 -3 26 5
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8783 0 0
2
5.90006e-315 5.32571e-315
0
7 Ground~
168 215 54 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3221 0 0
2
5.90006e-315 5.34643e-315
0
8 Op-Amp5~
219 292 144 0 5 11
0 5 3 7 6 4
0
0 0 64 0
5 LF353
12 -19 47 -11
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 589828
88 0 0 0 2 1 1 0
1 U
3215 0 0
2
5.90006e-315 5.3568e-315
0
9 Resistor~
219 298 67 0 2 5
0 3 4
0
0 0 864 0
2 2k
-7 -11 7 -3
2 RF
-6 -22 8 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7903 0 0
2
5.90006e-315 5.36716e-315
0
9 Resistor~
219 239 99 0 4 5
0 3 2 0 -1
0
0 0 864 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7121 0 0
2
5.90006e-315 5.37752e-315
0
9
1 0 3 0 0 8320 0 7 0 0 5 3
280 67
266 67
266 138
5 0 4 0 0 4096 0 6 0 0 7 2
310 144
341 144
1 1 5 0 0 12416 0 2 6 0 0 4
189 138
218 138
218 150
274 150
2 1 2 0 0 4224 0 8 5 0 0 4
239 81
239 41
215 41
215 48
1 2 3 0 0 0 0 8 6 0 0 3
239 117
239 138
274 138
1 2 2 0 0 0 0 1 2 0 0 3
206 159
206 148
189 148
2 0 4 0 0 8320 0 7 0 0 0 4
316 67
341 67
341 144
363 144
1 4 6 0 0 4224 0 3 6 0 0 2
292 169
292 157
1 3 7 0 0 4224 0 4 6 0 0 4
292 118
292 132
292 132
292 131
3
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
345 126 368 144
350 130 362 142
2 Vo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
280 84 307 108
285 88 301 104
2 +V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
280 179 307 203
285 183 301 199
2 -V
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1705266 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12401 0
4 1 10
1
335 144
0 2 0 0 3	0 10 0 0
1967280 8550464 100 100 0 0
77 66 767 156
0 322 800 570
767 66
77 66
767 66
767 156
0 0
0 0 0 0 0 0
12385 0
4 1e-06 10
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
