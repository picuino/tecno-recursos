��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  ��    S2      �  �� ��     S1      �  ����    L2      �  �Y�g    L1      �  � a � o     S1      �  � y � �     L1      �  )y 9�     L2                    ���  CBattery��  CValue  � �     9V         "@      �? V �� 	 CTerminal  �( �)              "@          �  �( �)                             � �4         ��      �� 	 CRailThru�  �( )       e       "@          �  �( 	)              "@            �$ ,          ����    ��  �H I        d                   �  �H 	I                             �D L          ����    ��  �� �       d        �          �  �� 	�                             �� �          ����    ��  CSPDT��  CToggle  ��(      "   �  �� ��                �          �  �� ��                �          �  � �                            �� �    %      ��    ��  �()      d                   �  �(	)                            �$,     )    ����    ��  �       d        �          �  � 	                            ��      ,    ����    ��  �� �       d        �          �  �� 	�                             �� �      /    ����    ��  �� �       d                   �  �� 	�                             �� �      2    ����    !�#�  �� ��       4   �  �� ��                �          �  �� ��                �          �  �� ��                             �| ��     6      ��    ��  �h i       d        �          �  �h 	i                             �d l      :    ����    ��  �HI      d        �          �  �H	I                            �DL     =    ����    ��  CBulb�  �H�I               �          �  �H�I     	          �            �<�T    A    ��      ��  �hi     	 d        �          �  �h	i     
                       �dl     D    ����    ��  ���      d        �          �  ��	�                            ���     G    ����    ?��  ����               �          �  ����               �            �|��    J    ��      ��  ���      d        �          �  ��	�                            ���     M    ����    ��   a 3 o     9V(          "@      �? V �  @ H A ]               "@
ףp=
��  �  @ t A �                 
ףp=
�?    4 \ L t      Q    ��      ?��  � ` � u               "@
ףp=
�?  �  � � � �                 
ףp=
��    � t � �      T  
 ��      ?��  ` u                 �          �  � �                             t $�      W    ��      !�#�  x @ � `      Y   �  h 0 } 1              "@
ףp=
�?  �  � 8 � 9              "@
ףp=
��  �  � ( � )                �            | $ � <      [     ��                  ���  CWire  �( �)       _�  �H �I        _�  �( �I         _�  �( �)        _�  �� ��       _�  �� ��        _�  �� ��       _�  �� ��       _�  �� �       _�  � �      _�  �(�)      _�  � �)       _�  � �      _�  �� ��       _�  �� ��        _�  �� ��       _�  �� ��       _�  �� ��        _�  �� ��       _�  �h �i       _�  �h ��        _�  �� ��       _�  �H�I      _�  �h�i     	 _�  �H�i      	 _�  �H�I     	 _�  ����      _�  ����       _�  ����      _�  ����      _�  @ 0 i 1       _�  @ 0 A I        _�  @ � A �        _�  @ � � �       _�  � � � �        _�  � � �       _�  � �        _�  � 8 � 9       _�  � 8 � a        _�  � ( )       _�  ( a                      �                              `  c  `      a      f        % % g & d & ' l ' j ) * *   i , - -   p / 0 0   o 2 3 3   6 6 r 7 u 7 8 m 8 s : ; ;   v = > >   A A v B y B w D E E   | G H H   J J } K z K } M N N   Q  Q R R � T � T U U � W � W X X � [ ~ [ \ \ � ] ] �   b  c a b  e & f d e  % h g i h , k ) l j k ' n 8 m o n 2 q / r p 6 q t : s u t 7 A = x D y w x B { K z | { G J M  [ ~ Q R � � � U � � � X � \ � � T ] � � W            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 