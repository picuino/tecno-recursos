��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  � i � w     S1      �  � i w     S2      �  Ya io     L1      �  �a	o    L1      �  ��	�    L2      �  � *�     S1      �  *'    S2                    ���  CBulb�� 	 CTerminal  HH I]                 �          �  Ht I�                              <\ Tt          ��      ��  CSPDT��  CToggle  � @ `          �  0 1                �          �  � ( � )              "@          �  � 8 � 9                             � $ <           ��    ��  x @ � `          �  h 0 } 1              "@          �  � 8 � 9                           �  � ( � )              "@            | $ � <            ��    ��  CBattery��  CValue   a 3 o     9V(          "@      �? V �  @ H A ]               "@          �  @ t A �                             4 \ L t      %    ��      �� 	 CRailThru�  0�E�      d                   �  4�I�               �            2�F�     )    ����    ��  �!�                          �  ����               �            ���    ,    ��      '��  0�E�      d        �          �  4�I�                            2�F�     /    ����    '��  0pEq      d        �          �  4pIq                            2lFt     2    ����    ��  P!Q               �          �  �P�Q               �            �D\    5    ��      '��  0PEQ      d        �          �  4PIQ                            2LFT     8    ����    '��  0p Eq       d        �          �  4p Iq                             2l Ft      ;    ����    ��  �� �       =   �  � �                �          �  �� ��                �          �  �� ��                             �� �     ?      ��    '��  0� E�       d                   �  4� I�                             2� F�      C    ����    '��  0� E�       d        �          �  4� I�                             2� F�      F    ����    '��  0E	      d        �          �  4I	                            2F     I    ����    '��  00E1      d                   �  40I1                            2,F4     L    ����    ��  �0      N   �                  �          �  �� ��      	          �          �  ��	                            ��     P      ��    '��  0� E�      	 d        �          �  4� I�      
                       2� F�      T    ����    '��  0P EQ       d                   �  4P IQ                             2L FT      W    ����    '��  00 E1       e       "@          �  40 I1              "@            2, F4      Z    ����    !�#�  � %     9V         "@      �? V �  �0 1              "@          �  �0 �1                            �$ �<     ^    ��                    ���  CWire  H0 II        a�  0 I1       a�  H� I�         a�  @ � I�        a�  @ � A �         a�  � ( � )       a�  � 8 � 9       a�  @ 0 A I        a�  @ 0 i 1       a�   �1�      a�  ��1�      a�  ����       a�  ����      a�  �P�Q      a�  �P�q       a�  �p1q      a�   P1Q      a�  �� ��       a�  �p ��        a�  �p 1q       a�  � )�       a�  (� )�        a�  (� 1�       a�  �� 1�       a�  �� ��        a�  �� ��       a�  ��	      a�  ��1       a�  �011      a�  (1	      a�  ( )	       a�   )      a�  �� 1�      	 a�  �� ��       	 a�  �� ��      	 a�  �0 �1       a�  �0 �Q        a�  �P 1Q       a�  0 11                     �                             b    d   c  g   h   j    h     g % i % & & f k ) * *   , , k - n - l / 0 0   q 2 3 3   5 5 r 6 o 6 r 8 9 9   u ; < <   ? ? v @ s @ A { A y C D D   x F G G    I J J   ~ L M M   P P � Q � Q R | R � T U U   � W X X   � Z [ [   ^ ^ � _ � _ c   b  e f d & e      j % i  , ) m / n l m - p 6 o q p 2 5 8 t @ u s t ; ? w v x w F z C { y z A } R | ~ } L � I �  P � � T � � � Q � _ � � � W ^ Z   "         �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 