��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  9aIo    L1      �  9�I�    L2      �  Y� j�     S1      �  Yj'    S2      �  � Y � g     S1      �  )I 9W     L1      �  )� 9�     L2      �  �I �W     S2                    ��� 	 CRailThru�� 	 CTerminal  p���      d                   �  t���               �            r���         ����    ��  CBulb�  L�a�                          �   �5�               �            4�L�        ��      ��  p���      d        �          �  t���                            r���         ����    ��  pp�q      d        �          �  tp�q                            rl�t         ����    ��  LPaQ               �          �   P5Q               �            4DL\    !    ��      ��  pP�Q      d        �          �  tP�Q                            rL�T     $    ����    ��  pp �q       d        �          �  tp �q                             rl �t      '    ����    ��  CSPDT��  CToggle  (� H�       *   �  D� Y�                �          �  � -�                �          �  � -�                             ,� D�     -      ��    ��  p� ��       d                   �  t� ��                             r� ��      1    ����    ��  p� ��       d        �          �  t� ��                             r� ��      4    ����    ��  p�	      d        �          �  t�	                            r�     7    ����    ��  p0�1      d                   �  t0�1                            r,�4     :    ����    )�+�  (H0      <   �  D Y               �          �  � -�      	          �          �  -	                            ,� D    >      ��    ��  p� ��      	 d        �          �  t� ��      
                       r� ��      B    ����    ��  pP �Q        d                   �  tP �Q                             rL �T      E    ����    ��  p0 �1       e       "@          �  t0 �1              "@            r, �4      H    ����    ��  CBattery��  CValue   D%     9V         "@      �? V �  <0 Q1              "@          �  0 %1                             $$ <<     N    ��      J�L�  3 q [      9V(          "@      �? V �  h X i m               "@          �  h � i �                �            \ l t �      R    ��      ��  CSPST+�  � 8 � X       U   �  � 0 � 1              "@          �  � 0 � 1                �            � , � 4      W      ��    ��  0 E                 �          �  \ q                �            D $\      Z    ��      ��  p �        	        �          �  � �                �            � $�      ]    ��      T�+�  �@ �`       _   �  x\ yq                �          �  x0 yE                 �            tD |\     a      ��                  ���  CWire  `�q�      d�   �q�      d�   ��       d�   �!�      d�   P!Q      d�   Pq       d�   pqq      d�  `PqQ      d�   � �       d�   p �        d�   p qq       d�  X� i�       d�  h� i�        d�  h� q�       d�   � q�       d�   � �        d�   � �       d�   	      d�   1       d�   0q1      d�  hq	      d�  h i	       d�  X i      d�   � q�      	 d�   � �       	 d�   � �      	 d�   0 1        d�   0 Q         d�   P qQ        d�  P0 q1       d�  h 0 i Y        d�  h 0 � 1       d�  � 0 1       d�  h � i �        d�  h � �       d�  p yq       d�  0 y1                     �                            e        e  h  f      k      ! ! l " i " l $ % %   o ' ( (   - - p . m . / u / s 1 2 2   r 4 5 5   y 7 8 8   x : ; ;   > > { ? ~ ? @ v @ | B C C   � E F F   � H I I   N N � O  O R � R S S � W � W X X � Z � Z [ [ � ] [ ] ^ ^ � a a � b � b   g  h f g  j " i k j  ! $ n . o m n ' - q p r q 4 t 1 u s t / w @ v x w : z 7 { y > z } B | ~ } ? � O  � � E N H � R � W X � S � � ^ ] a Z b   K         �%s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 