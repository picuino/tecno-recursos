CircuitMaker Text
5.6
Probes: 2
Vo
Transient Analysis
0 278 116 8421376
Vi_1
Transient Analysis
1 120 125 4227327
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 361
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1446 465
9961490 0
0
6 Title:
5 Name:
0
0
0
10
11 Signal Gen~
195 71 129 0 64 64
0 5 2 1 86 -10 10 9 0 0
0 0 0 0 0 0 0 1120403455 -1090519040 1056964608
0 0 0 1000593163 1008981771 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 100 -0.5 0.5 0 0 0 0.005 0.01 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -500m/500mV
-39 -31 38 -23
2 Vi
-7 -40 7 -32
0
0
44 %D %1 %2 DC 0 PULSE(-500m 500m 0 0 0 5m 10m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3277 0 0
2
44517.5 7
0
8 Op-Amp5~
219 239 130 0 5 11
0 2 4 6 7 3
0
0 0 80 0
5 LF353
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 0 2 1 1 0
1 U
4212 0 0
2
44517.5 6
0
7 Ground~
168 107 196 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4720 0 0
2
44517.5 5
0
2 +V
167 239 176 0 1 3
0 7
0
0 0 53616 180
4 -15V
-14 -1 14 7
3 Vi3
-10 0 11 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5551 0 0
2
44517.5 4
0
2 +V
167 239 101 0 1 3
0 6
0
0 0 53616 0
3 15V
-10 -14 11 -6
3 Vi4
-10 -24 11 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6986 0 0
2
44517.5 3
0
11 Terminal:A~
194 286 130 0 1 3
0 3
0
0 0 57584 180
2 Vo
-7 -13 7 -5
2 J1
-7 -23 7 -15
0
3 Vo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
8745 0 0
2
44517.5 2
0
10 Capacitor~
219 237 74 0 2 5
0 4 3
0
0 0 848 0
6 0.01uF
-22 -18 20 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9592 0 0
2
44517.5 1
0
7 Ground~
168 196 198 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8748 0 0
2
44517.5 0
0
9 Resistor~
219 146 124 0 2 5
0 5 4
0
0 0 880 0
4 100k
-13 -14 15 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
44517.5 10
0
9 Resistor~
219 239 35 0 2 5
0 4 3
0
0 0 880 0
4 1meg
-13 -14 15 -6
2 Rf
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
631 0 0
2
44517.5 8
0
11
2 0 3 0 0 4096 0 7 0 0 4 2
246 74
280 74
1 0 4 0 0 4096 0 7 0 0 5 2
228 74
197 74
2 0 4 0 0 0 0 2 0 0 5 2
221 124
197 124
2 1 3 0 0 8336 0 10 6 0 0 3
257 35
280 35
280 130
1 2 4 0 0 8320 0 10 9 0 0 4
221 35
197 35
197 124
164 124
1 1 2 0 0 8320 0 2 8 0 0 3
221 136
196 136
196 192
1 1 5 0 0 4224 0 9 1 0 0 2
128 124
102 124
5 1 3 0 0 0 0 2 6 0 0 2
257 130
280 130
3 1 6 0 0 4224 0 2 5 0 0 4
239 117
239 109
239 109
239 110
1 4 7 0 0 4224 0 4 2 0 0 2
239 161
239 143
2 1 2 0 0 0 0 1 3 0 0 3
102 134
107 134
107 190
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0.0401 0.06 0.0002 0.0002
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
2425688 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 10
0
2491180 8550464 100 100 0 0
77 66 767 156
0 322 800 570
472 66
77 66
767 66
767 156
0 0
0 0 0 0 0 0
12401 0
4 0.01 10
2
116 108
0 7 0 0 1	0 12 0 0
272 114
0 3 0 0 1	0 12 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
