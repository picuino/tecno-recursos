��  CCircuit��  CSerializeHack           ��  CPart  0   0       ���  CBattery��  CValue   !; /    9V(          "@      �? V �� 	 CTerminal  H I         U���!@�d��eݿ  �  H 4I I         ���A�(�d��e�?    < T 4         ��      ��  CDPDT��  CToggle  � H� h         �  x �        U���!@�d��e�?  �  x 8� 9          ���A�(�d��eݿ  �  � @� A       U���!@          �  � 0� 1          ���A�(�d��e�?  �  �  � !          ���A�          �  � �        U���!@�d��eݿ    � � D           �� ,   ��  CMotorEM�          U���!@(�d��e�?  �  4I          ���A�(�d��eݿ  �� 	 CMechTermc�p@^�����AtZ���      �<                  !     	 c�p@^���      �<    4        ��      bK�6�>c�p@^����{v���"3��5�c�p@^����{v�����  CBulb�  �	�              "@
ףp=
�?  �  �	�     	          �
ףp=
��    � ��     !  
 ��      ��  � �� �      
          �          �  � �� �     	          �            � �� �     $    ��      ��  CSPDT�  � �� �      '   �  p �� �             "@
ףp=
�?  �  � �� �     
          �          �  � �� �             "@
ףp=
��    � �� �     )      ��    �
�   �; �    9V(          "@      �? V �  H �I �              "@
ףp=
��  �  H �I �     	         �
ףp=
�?    < �T �     .    ��      �
�   � ; �     9V(          "@      �? V �  H � I �               "@          �  H � I �                             < � T �      2    ��      ��  � � � �                 �          �  � � � �                              � � � �      5    ��      ��  CSPST�  � ( � H       8   �  p   � !              "@          �  �   � !                �            �  � $      :      ��    ��  � 0 � E                 �          �  � \ � q                             � D � \      =    ��      �
�   I ; W     9V(          "@      �? V �  H 0 I E               "@          �  H \ I q                            < D T \      A    ��      �� 	 CPushMake��  CKey  � � � �       D   �  p � � �              "@          �  � � � �                �            � � � �      G      ��    ��  �  � 5              "@
ףp=
�?  �  � L� a                
ףp=
��    � 4� L     J  
 ��      �
�   9; G    9V(          "@      �? V �  H  I 5              "@
ףp=
��  �  H LI a               
ףp=
�?    < 4T L     N    ��      �� 
 CPushBreakE�  � � 6      Q   �  p �              "@
ףp=
�?  �  � �              "@
ףp=
��    � �      S      ��      0   0       ���  CWire  H y 	      V�  x y        V�  x 8y I       V�  H Hy I      V�  �  � !      V�  �  � 1       V�  � 0� 1      V�  � �        V�  � � A       V�  � � 	      V�  � 	      V��� 
 CCrossOver  � <� D        � @� A      V�c�  � <� D        � 0� I       V�  � HI      V�  H �� �     	 V�  � �	�     	 V�  �	�       V�  � �	�      V�  � �� �     
 V�  H �q �      V�  H �I �       V�  H � � �        V�  �   � !       V�  �   � 1        V�  H p � q       V�  H   I 1        V�  H   q !       V�  � � � �       V�  � � � �        V�  H � q �       V�  H � I �        V�  H `� a      V�  � �       V�  � � !       V�  H q       V�  H I !         0   0       �  0   0         0   0        W    Z  X   Y    b   ]   [   ^  a    g     ! j ! " " i $ l $ % % i ) m ) * * l + + k . n . / / h 2 x 2 3 3 o 5 v 5 6 6 o : t : ; ; p = q = > > r A s A B B r G w G H H u J { J K K y N } N O O y S | S T T z  X W   Z  Y  \ [ e  \ `  a b ^ _ `  b f  _ e d ] g e  / % h " k ! + j * $ n ) m . 3 6 ; q p = B > t A s : H v u 5 x G w 2 O K T { z J } S | N   0        �5s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 