��  CCircuit��  CSerializeHack           ��  CPart�� 	 CGroupBox  D�T�             �  $ ��             �  D$ T�              �  $ $ �                            ���  CBattery��  CDummyValue  �8�8    1.5V            �?      �? V �� 	 CTerminal  �(�=         �U  �?x����  �  ����     
  l�����   C�{z<    �<��         ��   �  ��  x8x8    1.5V            �?      �? V �  x(y=         eC  @          �  x�y�        �U  �?x���=    h<��         ��   �  �� 	 CFilament�  ��    1W            �?      �? W �  ��       k�����mN�VՂ<  �  )     
  l�����mN�VՂ�    ��(           ��`   �� 	 CPushMake��  CKey  �"�        �  �	        eC  @          �  �       k�����            ��!�     !    ����    ��  HH    1W            �?      �? W �  8M     	          �          �  ��               �            L��(     %      ��`   �� 
 CBattery9V�  � H� H    9V            "@      �? V �  � 8� M                �          �  ` 8a M              "@            L L� �     *    ��   �  ��  � �� �      ,  �  � ��              "@          �  � ��      	          �            � �� �     .    ����    �� 
 CVResistor��  CSlider  �i o�    	 �  �� ��     70            Y@ffffff�?    4 �  �� ��        8�W���!@,���
�?  �  t� ��         zd׾� �?,���
��    �� t�      5      ���   '��  �� ��     9V            "@      �? V �  �� ��              _���.���
�?  �  x� y�         8�W���!@3���
��    d� �h     9    ��   �  ��  �� ��     1W            �?      �? W �  �� ��         zd׾� �?.���
�?  �  � )�             _���.���
��    �N �      =      ��`   '��  � � � �     9V            "@      �? V �  � � � �                            �  X � Y �               "@            D � � h     A    ��   �  ��  CSPST��  CToggle  � @  d       D  �  � � � �              "@          �  � � � �                �            � b  �      G    ����P    ��  H� H�     1W            �?      �? W �  8� M�                �          �  �� ��                              LN ��      K      ��`                 ���  CWire  ()�      
 N�  ��)�     
 N�  x	      N�  xy)       N�  �      N�  �(�)      N�  �(��       N�  x���      N�  � 8�9      N�  ��9       N�  ` a 9       N�  ` �       N�  � 9     	 N�  � � ��        N�  X � � �       N�  �� ��       N�  (� )�        N�  �� )�       N�  x� y�        N�  x� ��       N�  �� ��         N�  � � 9�       N�  X � Y �                      �                             T    P  R    V  S    O ! ! Q " " S % [ % & & X * W * + Y + . . Z / / [ 5 b 5 6 6 ^ 9 ` 9 : a : = ^ = > > _ A \ A B e B G G ] H H d K d K L L c  P  O R ! Q  "  U  T V  U * X & W Z + Y . / % A c e G 6 = > ` 9 _ b : a 5 L \ H K ] B   ?         �4s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 