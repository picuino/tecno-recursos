CircuitMaker Text
5.6
Probes: 3
V1_1
Transient Analysis
0 89 86 4227327
V2_1
Transient Analysis
1 122 73 12615808
U1A_1
Transient Analysis
2 181 80 8421376
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1278 361
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 2 0.500000 0.500000
344 176 1446 465
9961490 0
0
6 Title:
5 Name:
0
0
0
6
7 Ground~
168 98 113 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9323 0 0
2
44525.2 5
0
11 Signal Gen~
195 48 90 0 64 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1092616192
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 1000 0 10 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -10/10V
-25 -30 24 -22
2 V1
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 10 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
317 0 0
2
44525.2 4
0
8 Op-Amp5~
219 155 79 0 5 11
0 4 3 6 7 5
0
0 0 80 0
5 LF353
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 0 2 1 1 0
1 U
3108 0 0
2
44525.2 3
0
2 +V
167 155 125 0 1 3
0 7
0
0 0 53360 180
4 -15V
-14 -1 14 7
3 Vi3
-10 0 11 8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4299 0 0
2
44525.2 2
0
2 +V
167 155 41 0 1 3
0 6
0
0 0 53360 0
3 15V
-10 -14 11 -6
3 Vi4
-10 -24 11 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9672 0 0
2
44525.2 1
0
2 +V
167 105 33 0 1 3
0 3
0
0 0 54128 0
2 5V
-8 -14 6 -6
2 V2
-8 -24 6 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7876 0 0
2
44525.2 0
0
6
1 2 3 0 0 8336 0 6 3 0 0 3
105 42
105 73
137 73
1 1 4 0 0 4240 0 2 3 0 0 2
79 85
137 85
1 2 2 0 0 8336 0 1 2 0 0 3
98 107
98 95
79 95
5 0 5 0 0 4240 0 3 0 0 0 2
173 79
195 79
3 1 6 0 0 4240 0 3 5 0 0 2
155 66
155 50
1 4 7 0 0 4240 0 4 3 0 0 2
155 110
155 92
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
143 121 174 145
150 127 166 143
2 -V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
143 15 168 39
147 19 163 35
2 +V
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
181 60 202 78
185 64 197 76
2 Vo
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2425688 1210432 100 100 0 0
0 0 0 0
0 74 161 144
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 10
0
2491180 8550464 100 100 0 0
77 66 767 156
0 322 800 570
472 66
77 66
767 66
767 156
0 0
0 0 0 0 0 0
12401 0
4 0.01 10
2
116 108
0 7 0 0 1	0 7 0 0
272 114
0 3 0 0 1	0 7 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
