��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  � Q � _     S2      �  ��    S2      �  �� ��     S1      �  ����    L2      �  �Y�g    L1      �  � a � o     S1      �  � y � �     L1      �  )y 9�     L2                    ���  CSPST��  CToggle  � 0  P          �� 	 CTerminal  � ( � )                �          �  � ( )                �            � $ � ,            ��    ��  CBattery��  CValue  � �     9V         "@      �? V �  �( �)              "@          �  �( �)                             � �4         ��      �� 	 CRailThru�  �( )       e       "@          �  �( 	)              "@            �$ ,           ����    ��  �H I        d                   �  �H 	I                             �D L      #    ����    ��  �� �       d        �          �  �� 	�                             �� �      &    ����    ��  CSPDT�  ��(      )   �  �� ��                �          �  �� ��                �          �  � �                            �� �    +      ��    ��  �()      d                   �  �(	)                            �$,     /    ����    ��  �       d        �          �  � 	                            ��      2    ����    ��  �� �       d        �          �  �� 	�                             �� �      5    ����    ��  �� �       d                   �  �� 	�                             �� �      8    ����    (��  �� ��       :   �  �� ��                �          �  �� ��                �          �  �� ��                             �| ��     <      ��    ��  �h i       d        �          �  �h 	i                             �d l      @    ����    ��  �HI      d        �          �  �H	I                            �DL     C    ����    ��  CBulb�  �H�I               �          �  �H�I     	          �            �<�T    G    ��      ��  �hi     	 d        �          �  �h	i     
                       �dl     J    ����    ��  ���      d        �          �  ��	�                            ���     M    ����    E��  ����               �          �  ����               �            �|��    P    ��      ��  ���      d        �          �  ��	�                            ���     S    ����    ��   a 3 o     9V(          "@      �? V �  @ H A ]               "@
ףp=
��  �  @ t A �                 
ףp=
�?    4 \ L t      W    ��      E��  � ` � u               "@
ףp=
�?  �  � � � �                 
ףp=
��    � t � �      Z  
 ��      E��  ` u                 �          �  � �                             t $�      ]    ��      (��  x @ � `      _   �  h 0 } 1              "@
ףp=
�?  �  � 8 � 9              "@
ףp=
��  �  � ( � )                �            | $ � <      a     ��                  ���  CWire  � ( � )       e�  ( a        e�  ( )       e�  �( �)       e�  �H �I        e�  �( �I         e�  �( �)        e�  �� ��       e�  �� ��        e�  �� ��       e�  �� ��       e�  �� �       e�  � �      e�  �(�)      e�  � �)       e�  � �      e�  �� ��       e�  �� ��        e�  �� ��       e�  �� ��       e�  �� ��        e�  �� ��       e�  �h �i       e�  �h ��        e�  �� ��       e�  �H�I      e�  �h�i     	 e�  �H�i      	 e�  �H�I     	 e�  ����      e�  ����       e�  ����      e�  ����      e�  @ 0 i 1       e�  @ 0 A I        e�  @ � A �        e�  @ � � �       e�  � � � �        e�  � � �       e�  � �        e�  � 8 � 9       e�  � 8 � a                      �                             f    h   i  l  i   ! !   j # $ $   o & ' '   + + p , m , - u - s / 0 0   r 2 3 3   y 5 6 6   x 8 9 9   < < { = ~ = > v > | @ A A    C D D   G G  H � H � J K K   � M N N   P P � Q � Q � S T T   W � W X X � Z � Z [ [ � ] g ] ^ ^ � a � a b b � c c f c  h ]  g    k # l j k  n , o m n & + q p r q 2 t / u s t - w > v x w 8 z 5 { y < z } @ | ~ } = G C � J � � � H � Q � � � M P S � a � W X � � � [ � � � ^ � b � � Z            �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 