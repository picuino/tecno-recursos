CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
21 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1278 659
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
37 C:\Archivos de programa\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
10
8 Op-Amp5~
219 317 149 0 5 11
0 5 3 8 7 3
0
0 0 64 0
5 UA741
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
3409 0 0
2
5.89937e-315 5.26354e-315
0
10 Capacitor~
219 233 155 0 2 5
0 5 4
0
0 0 576 180
6 0.01uF
-21 -18 21 -10
2 C2
-7 -19 7 -11
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3951 0 0
2
5.89937e-315 5.30499e-315
0
11 Signal Gen~
195 105 160 0 64 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162722
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 64 0
5 -1/1V
-18 -30 17 -22
2 Vi
-6 -31 8 -23
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 1 0 0
1 V
8885 0 0
2
5.89937e-315 5.32571e-315
0
7 Ground~
168 276 220 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3780 0 0
2
5.89937e-315 5.34643e-315
0
7 Ground~
168 136 220 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9265 0 0
2
5.89937e-315 5.3568e-315
0
2 +V
167 317 118 0 1 3
0 8
0
0 0 53344 0
3 15V
-9 -25 12 -17
2 V1
-6 -14 8 -6
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9442 0 0
2
5.89937e-315 5.36716e-315
0
2 +V
167 317 186 0 1 3
0 7
0
0 0 53344 180
4 -15V
-12 10 16 18
2 V2
-6 -1 8 7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9424 0 0
2
5.89937e-315 5.37752e-315
0
10 Capacitor~
219 166 155 0 2 5
0 6 4
0
0 0 576 0
6 0.01uF
-22 -18 20 -10
2 C1
-7 -20 7 -12
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9968 0 0
2
5.89937e-315 5.38788e-315
0
9 Resistor~
219 276 187 0 3 5
0 2 5 -1
0
0 0 608 90
5 22.5k
11 0 46 8
2 R1
4 -3 18 5
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9281 0 0
2
5.89937e-315 5.39306e-315
0
9 Resistor~
219 241 68 0 2 5
0 4 3
0
0 0 608 0
6 11.25k
-21 -14 21 -6
2 R2
-7 -12 7 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8464 0 0
2
5.89937e-315 5.40342e-315
0
11
2 0 3 0 0 12288 0 1 0 0 2 4
299 143
276 143
276 91
375 91
2 5 3 0 0 8336 0 10 1 0 0 4
259 68
375 68
375 149
335 149
1 0 4 0 0 8320 0 10 0 0 7 3
223 68
195 68
195 155
1 1 2 0 0 4096 0 9 4 0 0 4
276 205
276 215
276 215
276 214
2 0 5 0 0 4096 0 9 0 0 6 2
276 169
276 155
1 1 5 0 0 4224 0 2 1 0 0 2
242 155
299 155
2 2 4 0 0 0 0 2 8 0 0 2
224 155
175 155
1 1 6 0 0 4224 0 8 3 0 0 2
157 155
136 155
1 4 7 0 0 4224 0 7 1 0 0 2
317 171
317 162
1 3 8 0 0 4224 0 6 1 0 0 2
317 127
317 136
1 2 2 0 0 4224 0 5 3 0 0 2
136 214
136 165
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
91 118 118 142
96 122 112 138
2 Vi
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
299 93 336 117
309 101 325 117
2 +V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
298 174 335 198
308 182 324 198
2 -V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
346 122 383 146
356 130 372 146
2 Vo
0
9 0 0
0
0
2 V1
-0.7 -1.5 -0.02
0
0 0 0
100 0 10 10000
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
5768164 1210432 100 100 0 0
0 0 0 0
0 107 161 177
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 5e-06 10
0
5309400 4421696 100 100 0 0
77 66 779 156
-4 333 798 572
545 66
311 66
779 84
779 111
0 0
0 0 0 0 0 0
12403 0
4 500 1000
1
369 149
0 3 0 0 3	0 12 0 0
6030466 4421696 100 100 0 0
77 66 767 156
-4 333 798 572
86 66
77 66
767 97
767 97
0 0
0 0 0 0 0 0
12401 0
4 20 0.5
1
324 112
0 5 0 0 3	0 12 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
